netcdf vrc {

    dimensions:
        record = unlimited,
        z = 1,
	x = 125,
	y = 105,
        nav = 1,
        namelen = 132;
		
    variables:
        //	NOWRAD 2D radar

	float                                  
            ref(record,z,y,x);
            ref:navigation_dim = "nav";
            ref:record = "valtime, reftime";
            ref:_FillValue = 1.e+37f;
            ref:long_name="NOWRAD 2D radar reflectivity";
            ref:units="dBZ";
            ref:valid_range= -50.f, 100.f;
            ref:LAPS_var="REF";
            ref:lvl_coord="MSL";
	    ref:LAPS_units="DBZ";

        //      2D minimum radar distance

        float
            dis(record,z,y,x);
            dis:navigation_dim = "nav";
            dis:record = "valtime, reftime";
            dis:_FillValue = 1.e+37f;
            dis:long_name="NOWRAD 2D minimum radar distance";
            dis:units="dBZ";
            dis:valid_range= 0.f, 1000000.f;
            dis:LAPS_var="DIS";
            dis:lvl_coord="MSL";
            dis:LAPS_units="m";
                	        
        //	LAPS variables

        long
            imax,
            jmax,
            kmax,
            kdim;

        char
            ref_comment(record,z,namelen),
            dis_comment(record,z,namelen),
            asctime(record,namelen);

			
        //	inventory variables

        short
            ref_fcinv(record, z);
            ref_fcinv:_FillValue= 0s;
              	
        short
            dis_fcinv(record, z);
            dis_fcinv:_FillValue= 0s;
              	
        //	list of grid levels

        float 
            level(z);
            level:long_name="level of data";
	    level:units = "hectopascals";
                    	
        //      validtime of the grid 

        double
            valtime(record);
            valtime:long_name = "valid time";
            valtime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      reference time of the process

        double
            reftime(record);
            reftime:long_name = "reference time";
            reftime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      nice name for originating center

        char
            origin_name(namelen);

        //      nice name for process

        char
            process_name(namelen);

        //      nice name for grid description instance
        char
            grid_name(namelen);

        //      basic assumption about earth shape
        char
            earth_shape(namelen);

        // navigation variables using 
        // WMO FM 92-VIII Ext.GRIB specification names
  
        char    grid_type(nav, namelen);
                grid_type:long_name = "GRIB-1 grid type";
  
        char    x_dim(nav, namelen);
                x_dim:long_name = "longitude dimension";
  
        char    y_dim(nav, namelen);
                y_dim:long_name = "latitude dimension";
  
        short   Nx(nav);
                Nx:long_name = "number of x points";
  
        short   Ny(nav);
                Ny:long_name =  "number of y points";
  
        float   La1(nav);
                La1:long_name = "first latitude";
                La1:units = "degrees_north";
  
        float   Lo1(nav);
                Lo1:long_name = "first longitude";
                Lo1:units = "degrees_east" ;
    
        float   LoV(nav);
                LoV:long_name = "orientation of grid" ;
                LoV:units = "degrees_east";
  
        float   Latin1(nav);
                Latin1:long_name = "orientation of grid" ;
                Latin1:units = "degrees_north";

        float   Latin2(nav);
                Latin2:long_name = "orientation of grid" ;
                Latin2:units = "degrees_north";

        float   Dx(nav);
                Dx:long_name = "x grid increment";
                Dx:units = "kilometers";
  
        float   Dy(nav);
                Dy:long_name = "y grid increment";
                Dy:units = "kilometers";
  
        // end of navigation variables

        :Conventions = "NUWG";
        :history = "created by LAPS Branch of FSL";
        :record = "valtime, reftime";
        :title = "LAPS vrc file - NOWRAD 2D radar";
        :version = 3;

    data:

        earth_shape     = "spherical radius";
        grid_name       = "LAPS vrc file - NOWRAD 2D radar";
        process_name    = "LAPS - Local Analysis and Prediction System";
        x_dim           = "x";
        y_dim           = "y";
}                       
