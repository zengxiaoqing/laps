// ---------------------------------------------------------------------------
// This software is in the public domain, furnished "as is", without technical
// support, and with no warranty, express or implied, as to its usefulness for
// any purpose.
//
// laps.cdl  	Local Analysis and Prediction System Model
//
// Author: Tom Kent + Jim Ramer
// ---------------------------------------------------------------------------
//
// A few notes about this cdl file:
//
// - The navigation info is not used right now. It probably will be in the
//   future and will be updated at that time.
//
// - "enumField" attribute has been eliminated.  To account for this,
//   a new DataField table exists within the GridKeyServer.
//   
// - The "enumLevelType" attribute has been eliminated.  Also, there is no
//   longer a separate netCDF variable for each level type that a given
//   physical parameter is available for.  To account for this, each variable
//   will be accompanied by a metadata variable that will contain a list
//   of levels that this variable is available for, encoded as character
//   data.  The accessor code has been updated to decode and cache this the
//   the first time it encounters a netCDF file from a given source.
//   All known grid level types are now registered in the DataGridLevel
//   table within the GridKeyServer.
//
// - For each physical parameter represented here, there is two pieces of
//   metadata meant to describe which levels it is available on.  The
//   attribute `levels' is meant to be a human readable format that someone
//   doing a ncdump can see.  The variable `xxxLevels' is the data that
//   is parsed by the accessor to determine which 2d slab corresponds to
//   which level.
//
// - The _n3D attribute is how many 2d slabs should be read in to get a
//   three-dimensional description of this variable.  This will be used
//   later to optimize access for cross sections and soundings.
//
// - The inventory variable is 2d based on record (valid time) and
//   level.  There is a separate inventory variable for each
//   meteorological variable.
// 
// - The forecast times are stored in the variable valtimeMINUSreftime,
//   which is dimensioned n_valtimes in size.  n_valtimes should
//   correspond to the number of records in a completely full file.
//
// - The units and valid ranges are being checked for accuracy and will be
//   updated soon if need be. 
//

netcdf laps
    {

    dimensions:
	record 		= UNLIMITED;
	n_valtimes	= 1;
	data_variables 	= 46;
	namelen	 	= 132;
	charsPerLevel 	= 10;
	x = 199,
	y = 247,

        // arbitrary counters for number of levels
        levels_1	= 1;
        levels_2	= 2;
        levels_3	= 3;
        levels_21	= 21;
        levels_22	= 22;


    variables:
        
	//      Geopotential height
	float
	    gh(record, levels_21, y, x);
	    gh:long_name = "Geopotential height";
	    gh:units = "geopotential meters";
	    gh:valid_range = 0.f, 10000.f;
	    gh:_FillValue = -99999.f;
	    gh:_n3D = 21;
            gh:levels = "MB 1100-100 by 50";
        char
            ghLevels(levels_21, charsPerLevel);
        char
            ghInventory(n_valtimes, levels_21);
	    

	//	Relative Humidity	
	float
	    rh(record, levels_22, y, x);
	    rh:long_name = "Relative Humidity";
	    rh:units = "percent";
	    rh:valid_range = 0.f, 100.f;
	    rh:_FillValue = -99999.f;
	    rh:_n3D = 22;
            rh:levels = "SFC  MB 1100-100 by 50";
        char
            rhLevels(levels_22, charsPerLevel);
        char
            rhInventory(n_valtimes, levels_22);    


	//	Temperature 	
  	float
	    t(record, levels_22, y, x);
	    t:long_name = "Temperature";
	    t:units = "degrees K";
	    t:valid_range = 0.f, 400.f;
	    t:_FillValue = -99999.f;
	    t:_n3D = 22;
            t:levels = "SFC  MB 1100-100 by 50";
        char
            tLevels(levels_22, charsPerLevel);
        char
            tInventory(n_valtimes, levels_22);


	//	u wind component
	float
	    uw(record, levels_22, y, x);
	    uw:long_name = "u wind component";
	    uw:units = "meters/second";
	    uw:valid_range = -300.f, 300.f;
	    uw:_FillValue = -99999.f;
	    uw:_n3D = 22;
            uw:levels = "SFC  MB 1100-100 by 50";
        char
            uwLevels(levels_22, charsPerLevel);
        char
            uwInventory(n_valtimes, levels_22);

	
	//	v wind component
	float
	    vw(record, levels_22, y, x);
	    vw:long_name = "v wind component";
	    vw:units = "meters/second";
	    vw:valid_range = -300.f, 300.f;
	    vw:_FillValue = -99999.f;
	    vw:_n3D = 22;
            vw:levels = "SFC  MB 1100-100 by 50";
        char
            vwLevels(levels_22, charsPerLevel);
        char
            vwInventory(n_valtimes, levels_22);

	
	//	pressure vertical velocity 
	float
	    pvv(record, levels_22, y, x);
	    pvv:long_name = "Pressure vertical velocity";
	    pvv:units = "Pa/s";
	    pvv:valid_range = -10.f, 10.f;
	    pvv:_FillValue = -99999.f;
	    pvv:_n3D = 22;
            pvv:levels = "SFC  MB 1100-100 by 50";
        char
            pvvLevels(levels_22, charsPerLevel);
        char
            pvvInventory(n_valtimes, levels_22);
	

        //      specific humidity
        float
            sh(record,levels_21,y,x);
            sh:long_name="specific humidity";
            sh:units="kg/kg";
            sh:valid_range= 0.f, 0.1000f;
            sh:_FillValue = -99999.f;
	    sh:_n3D = 21;
            sh:levels = "MB 1100-100 by 50";
        char
            shLevels(levels_21, charsPerLevel);
        char
            shInventory(n_valtimes, levels_21);


        //      LAPS radar reflectivity 
        float
            rr(record,levels_21,y,x);
            rr:long_name="LAPS radar reflectivity";
            rr:units="dBZ";
            rr:valid_range= -200.f, 200.f;
            rr:_FillValue = -99999.f;
	    rr:_n3D = 21;
            rr:levels = "MB 1100-100 by 50";
        char
            rrLevels(levels_21, charsPerLevel);
        char
            rrInventory(n_valtimes, levels_21);

        
        //      precipitation type
        float
            ptyp(record,levels_21,y,x);
            ptyp:long_name="precipitation type";
            ptyp:units="none";
            ptyp:valid_range= -200.f, 200.f;
            ptyp:_FillValue = -99999.f;
	    ptyp:_n3D = 21;
            ptyp:levels = "MB 1100-100 by 50";
        char
            ptypLevels(levels_21, charsPerLevel);
        char
            ptypInventory(n_valtimes, levels_21);

        
        //      cloud type
        float
            ctyp(record,levels_21,y,x);
            ctyp:long_name="cloud type";
            ctyp:units="none";
            ctyp:valid_range= -200.f, 200.f;
            ctyp:_FillValue = -99999.f;
	    ctyp:_n3D = 21;
            ctyp:levels = "MB 1100-100 by 50";
        char
            ctypLevels(levels_21, charsPerLevel);
        char
            ctypInventory(n_valtimes, levels_21);


        //      fractional cloud cover pressure coord
        float
            ccpc(record,levels_21,y,x);
            ccpc:long_name="fractional cloud cover pressure coord";
            ccpc:units="fractional";
            ccpc:valid_range= 0.f, 100.f;
            ccpc:_FillValue = -99999.f;
	    ccpc:_n3D = 21;
            ccpc:levels = "MB 1100-100 by 50";
        char
            ccpcLevels(levels_21, charsPerLevel);
        char
            ccpcInventory(n_valtimes, levels_21);
        
        
        //      cloud liquid water
        float
            cw(record,levels_21,y,x);
            cw:long_name="cloud liquid water";
            cw:units="grams/meter**3";
            cw:valid_range= 0.f, 100.f;
            cw:_FillValue = -99999.f;
	    cw:_n3D = 21;
            cw:levels = "MB 1100-100 by 50";
        char
            cwLevels(levels_21, charsPerLevel);
        char
            cwInventory(n_valtimes, levels_21);


        //      cloud ice
        float
            cice(record,levels_21,y,x);
            cice:long_name="cloud ice";
            cice:units="grams/meter**3";
            cice:valid_range= 0.f, 100.f;
            cice:_FillValue = -99999.f;
	    cice:_n3D = 21;
            cice:levels = "MB 1100-100 by 50";
        char
            ciceLevels(levels_21, charsPerLevel);
        char
            ciceInventory(n_valtimes, levels_21);
 
        
        //      hydrometeor concentration
        float
            hyc(record,levels_21,y,x);
            hyc:long_name="hydrometeor concentration";
            hyc:units="grams/meter**3";
            hyc:valid_range= 0.f, 100.f;
            hyc:_FillValue = -99999.f;
	    hyc:_n3D = 21;
            hyc:levels = "MB 1100-100 by 50";
        char
            hycLevels(levels_21, charsPerLevel);
        char
            hycInventory(n_valtimes, levels_21);


        //      Pressure         //
        float
            p(record,levels_2,y,x);
            p:long_name="pressure";
            p:units="pascals";
            p:valid_range= 0.f, 1000.f;
            p:_FillValue = -99999.f;
	    p:_n3D = 1;
            p:levels = "SFC  FH 1500";
        char
            pLevels(levels_2, charsPerLevel);
        char
            pInventory(n_valtimes, levels_2);


        //      MSL Pressure            // 
        float
            mslp(record,levels_1,y,x);
            mslp:long_name="Mean Sea Level Pressure";
            mslp:units="pascals";
            mslp:valid_range= -20000.f, 20000.f;
            mslp:_FillValue = -99999.f;
	    mslp:_n3D = 0;
            mslp:levels = "SFC";
        char
            mslpLevels(levels_1, charsPerLevel);
        char
            mslpInventory(n_valtimes, levels_1);

        
        //      surface dewpoint temperature    // 
        float
            dpt(record,levels_1,y,x);
            dpt:long_name="surface dewpoint temperature";
            dpt:units="degrees kelvin";
            dpt:valid_range= -75.f, 125.f;
            dpt:_FillValue = -99999.f;
	    dpt:_n3D = 0;
            dpt:levels = "SFC";
        char
            dptLevels(levels_1, charsPerLevel);
        char
            dptInventory(n_valtimes, levels_1);


        //     surface Potential temperature   // 
        float
            pot(record,levels_1,y,x);
            pot:long_name="potential temperature";
            pot:units="degrees Kelvin";
            pot:valid_range= -75.f, 125.f;
            pot:_FillValue = -99999.f;
	    pot:_n3D = 0;
            pot:levels = "SFC";
        char
            potLevels(levels_1, charsPerLevel);
        char
            potInventory(n_valtimes, levels_1);


        //      Cloud Ceiling           //
         float
            cc(record,levels_2,y,x);
            cc:long_name="cloud ceiling";
            cc:units="meters";
            cc:valid_range= -20000.f, 20000.f;
            cc:_FillValue = -99999.f;
	    cc:_n3D = 0;
            cc:levels = "SFC  MSL";
        char
            ccLevels(levels_2, charsPerLevel);
        char
            ccInventory(n_valtimes, levels_2);


        //      Temperature Advection   // 
        float
            tadv(record,levels_1,y,x);
            tadv:long_name="temperature advection";
            tadv:units="degrees Kelvin/second";
            tadv:valid_range= -20000.f, 20000.f;
            tadv:_FillValue = -99999.f;
	    tadv:_n3D = 0;
            tadv:levels = "SFC";
        char
            tadvLevels(levels_1, charsPerLevel);
        char
            tadvInventory(n_valtimes, levels_1);


        //      equivalent potential temperature  // 
        float
            ept(record,levels_1,y,x);
            ept:long_name="equivalent potential temperature";
            ept:units="degrees Kelvin";
            ept:valid_range= -20000.f, 20000.f;
            ept:_FillValue = -99999.f;
	    ept:_n3D = 0;
            ept:levels = "SFC";
        char
            eptLevels(levels_1, charsPerLevel);
        char
            eptInventory(n_valtimes, levels_1);


        //      integrated liquid water 
        float
            ilw(record,levels_1,y,x);
            ilw:long_name="integrated liquid water";
            ilw:units="grams/meter**2";
            ilw:valid_range= 0.f, 100.f;
            ilw:_FillValue = -99999.f;
	    ilw:_n3D = 0;
            ilw:levels = "SFC";
        char
            ilwLevels(levels_1, charsPerLevel);
        char
            ilwInventory(n_valtimes, levels_1);


        //      moisture convergence            // 
        float
            mcon(record,levels_1,y,x);
            mcon:long_name="moisture convergence";
            mcon:units="grams/kilogram/seconds";
            mcon:valid_range= -20000.f, 20000.f;
            mcon:_FillValue = -99999.f;
	    mcon:_n3D = 0;
            mcon:levels = "SFC";
        char
            mconLevels(levels_1, charsPerLevel);
        char
            mconInventory(n_valtimes, levels_1);


        //      potential temperature advection         // 
        float
            pta(record,levels_1,y,x);
            pta:long_name="potential temperature advection";
            pta:units="kilograms/second";
            pta:valid_range= -20000.f, 20000.f;
            pta:_FillValue = -99999.f;
	    pta:_n3D = 0;
            pta:levels = "SFC";
        char
            ptaLevels(levels_1, charsPerLevel);
        char
            ptaInventory(n_valtimes, levels_1);


        //      lifted index            // 
        float
            sli(record,levels_1,y,x);
            sli:long_name="lifted index";
            sli:units="degrees Kelvin";
            sli:valid_range= -20000.f, 20000.f;
            sli:_FillValue = -99999.f;
	    sli:_n3D = 0;
            sli:levels = "SFC";
        char
            sliLevels(levels_1, charsPerLevel);
        char
            sliInventory(n_valtimes, levels_1);

	
	//	Heat Index	  
        float 
            hidx(record, levels_1,y, x);
            hidx:long_name = "Heat index" ;
            hidx:units = "degrees Kelvin" ;
            hidx:valid_range = 0.f, 300.f;
            hidx:_FillValue = -99999.f;
	    hidx:_n3D = 0;
            hidx:levels = "SFC";
        char
            hidxLevels(levels_1, charsPerLevel);
        char
            hidxInventory(n_valtimes, levels_1);


        //      colorado severe storm index     //
        float
            cssi(record,levels_1,y,x);
            cssi:long_name="colorado severe storm index";
            cssi:units="          ";
            cssi:valid_range= -20000.f, 20000.f;
            cssi:_FillValue = -99999.f;
 	    cssi:_n3D = 0;
            cssi:levels = "SFC";
        char
            cssiLevels(levels_1, charsPerLevel);
        char
            cssiInventory(n_valtimes, levels_1);

 
        //      positive buoyant energy         //
        float
            pbe(record,levels_1,y,x);
            pbe:long_name="positive buoyant energy";
            pbe:units="joules/kilogram";
            pbe:valid_range= -20000.f, 20000.f;
            pbe:_FillValue = -99999.f;
 	    pbe:_n3D = 0;
            pbe:levels = "SFC";
        char
            pbeLevels(levels_1, charsPerLevel);
        char
            pbeInventory(n_valtimes, levels_1);


        //      negative buoyant energy         // 
         float
            nbe(record,levels_1,y,x);
            nbe:long_name="negative buoyant energy";
            nbe:units="joules/kilogram";
            nbe:valid_range= -20000.f, 20000.f;
            nbe:_FillValue = -99999.f;
 	    nbe:_n3D = 0;
            nbe:levels = "SFC";
        char
            nbeLevels(levels_1, charsPerLevel);
        char
            nbeInventory(n_valtimes, levels_1);


         //      visability              //
         float
            vis(record,levels_1,y,x);
            vis:long_name="visibility";
            vis:_FillValue = -99999.f;
            vis:units="meters";
            vis:valid_range= -20000.f, 20000.f;
 	    vis:_n3D = 0;
            vis:levels = "SFC";
        char
            visLevels(levels_1, charsPerLevel);
        char
            visInventory(n_valtimes, levels_1);


        //      LAPS cloud cover 
        float
            ccov(record,levels_1,y,x);
            ccov:long_name="LAPS cloud cover";
            ccov:units="none";
            ccov:valid_range= 0.f, 100.f;
            ccov:_FillValue = -99999.f;
 	    ccov:_n3D = 0;
            ccov:levels = "SFC";
        char
            ccovLevels(levels_1, charsPerLevel);
        char
            ccovInventory(n_valtimes, levels_1);

        
        //      cloud base 
        float
            cb(record,levels_1,y,x);
            cb:long_name="LAPS cloud base";
            cb:units="meters";
            cb:valid_range= -200.f, 200.f;
            cb:_FillValue = -99999.f;
 	    cb:_n3D = 0;
            cb:levels = "SFC";
        char
            cbLevels(levels_1, charsPerLevel);
        char
            cbInventory(n_valtimes, levels_1);


        //      cloud top 
        float
            ctop(record,levels_1,y,x);
            ctop:long_name="LAPS cloud top";
	    ctop:units="meters";
            ctop:valid_range= -200.f, 200.f;
            ctop:_FillValue = -99999.f;
 	    ctop:_n3D = 0;
            ctop:levels = "SFC";
        char
            ctopLevels(levels_1, charsPerLevel);
        char
            ctopInventory(n_valtimes, levels_1);


        //       Max echo tops 
        float
            mret(record,levels_1,y,x);
            mret:long_name="maximum radar echo tops";
            mret:units="meters";
            mret:valid_range= 0.f, 0.100f;
            mret:_FillValue = -99999.f;
 	    mret:_n3D = 0;
            mret:levels = "SFC";
        char
            mretLevels(levels_1, charsPerLevel);
        char
            mretInventory(n_valtimes, levels_1);


        //      Low Level Reflectivity 
        float
            llr(record,levels_1,y,x);
            llr:long_name="low level reflectivity";
            llr:units="dBZ";
            llr:valid_range= 0.f, 0.100f;
            llr:_FillValue = -99999.f;
 	    llr:_n3D = 0;
            llr:levels = "SFC";
        char
            llrLevels(levels_1, charsPerLevel);
        char
            llrInventory(n_valtimes, levels_1);
        
        
        //      helicity 
        float
            heli(record,levels_1,y,x);
            heli:long_name="helicity";
            heli:units="meters / second**2";
            heli:valid_range= 0.f, 0.100f;
            heli:_FillValue = -99999.f;
 	    heli:_n3D = 0;
            heli:levels = "SFC";
        char
            heliLevels(levels_1, charsPerLevel);
        char
            heliInventory(n_valtimes, levels_1);

        
        //      integrated total precip water 
        float
            tpw(record,levels_1,y,x);
            tpw:long_name="integrated total precipitable water";
            tpw:units="meters";
            tpw:valid_range= 0.f, 0.100f;
            tpw:_FillValue = -99999.f;
 	    tpw:_n3D = 0;
            tpw:levels = "SFC";
        char
            tpwLevels(levels_1, charsPerLevel);
        char
            tpwInventory(n_valtimes, levels_1);

        
        //      60 min snow accumulation 
        float
            s1hr(record,levels_1,y,x);
            s1hr:long_name="LAPS 60 minute snow accum.";
            s1hr:units="meters";
            s1hr:valid_range= -200.f, 200.f;
            s1hr:_FillValue = -99999.f;
 	    s1hr:_n3D = 0;
            s1hr:levels = "SFC";
        char
            s1hrLevels(levels_1, charsPerLevel);
        char
            s1hrInventory(n_valtimes, levels_1);

        
        //      storm total accumulation 
        float
            stot(record,levels_1,y,x);
            stot:long_name="storm total snow accumulation";
            stot:units="meters";
            stot:valid_range= -200.f, 200.f;
            stot:_FillValue = -99999.f;
 	    stot:_n3D = 0;
            stot:levels = "SFC";
        char
            stotLevels(levels_1, charsPerLevel);
        char
            stotInventory(n_valtimes, levels_1);

        
        //      60 minute precip accumulation 
        float
            pc(record,levels_1,y,x);
            pc:long_name="LAPS 60 minute precip. accum.";
            pc:units="meters";
            pc:valid_range= -200.f, 200.f;
            pc:_FillValue = -99999.f;
 	    pc:_n3D = 0;
            pc:levels = "SFC";
        char
            pcLevels(levels_1, charsPerLevel);
        char
            pcInventory(n_valtimes, levels_1);

        
        //      storm total precip accum 
        float
            stpa(record,levels_1,y,x);
            stpa:long_name="storm total precip. accum.";
            stpa:units="meters";
            stpa:valid_range= -200.f, 200.f;
            stpa:_FillValue = -99999.f;
 	    stpa:_n3D = 0;
            stpa:levels = "SFC";
        char
            stpaLevels(levels_1, charsPerLevel);
        char
            stpaInventory(n_valtimes, levels_1);


        //      LAPS surface precip type 
        float
            spt(record,levels_1,y,x);
            spt:long_name="LAPS precip type";
            spt:units="none";
            spt:valid_range= -200.f, 200.f;
            spt:_FillValue = -99999.f;
 	    spt:_n3D = 0;
            spt:levels = "SFC";
        char
            sptLevels(levels_1, charsPerLevel);
        char
            sptInventory(n_valtimes, levels_1);


        //   LAPS surface precip type - low level radar reflectivity modified 
        float
            ptt(record,levels_1,y,x);
            ptt:long_name="LAPS precip type - LL radar ref modified";
            ptt:units="none";
            ptt:valid_range= -200.f, 200.f;
            ptt:_FillValue = -99999.f;
 	    ptt:_n3D = 0;
            ptt:levels = "SFC";
        char
            pttLevels(levels_1, charsPerLevel);
        char
            pttInventory(n_valtimes, levels_1);


        //  	Fire Index 
        float
            fd(record,levels_1,y,x);
            fd:long_name="Fire Index";
            fd:units="none";
            fd:valid_range= 0.f, 20.f;
            fd:_FillValue = -99999.f;
 	    fd:_n3D = 0;
            fd:levels = "SFC";
        char
            fdLevels(levels_1, charsPerLevel);
        char
            fdInventory(n_valtimes, levels_1);

       
        //     snow cover 
        float
            scp(record,levels_1,y,x);
            scp:long_name="snow cover percentage";
            scp:units="none";
            scp:valid_range= 0.f, 1.0f;
            scp:_FillValue = -99999.f;
 	    scp:_n3D = 0;
            scp:levels = "SFC";
        char
            scpLevels(levels_1, charsPerLevel);
        char
            scpInventory(n_valtimes, levels_1);


        //      soil moisture 
        float
            smc(record,levels_3,y,x);
            smc:long_name="soil moisture";
            smc:units="meter/meter";
            smc:valid_range= -200.f, 200.f;
            smc:_FillValue = -99999.f;
 	    smc:_n3D = 0;
            smc:levels = "BLS 1 2 3";
        char
            smcLevels(levels_3, charsPerLevel);
        char
            smcInventory(n_valtimes, levels_3);


	//	forecast times
        int
            valtimeMINUSreftime(n_valtimes);
            valtimeMINUSreftime:units = "seconds";

	//	time the data is valid at
	double	
	    valtime(record);
	    valtime:long_name = "valid time";
	    valtime:units = "seconds since (1970-1-1 00:00:00.0)";

	
	//	reference time of the model
	double	
	    reftime(record);
	    reftime:long_name = "reference time";
	    reftime:units = "seconds since (1970-1-1 00:00:00.0)";

	
	//	nice name for originating center
	char
	    origin(namelen);

	
	//	nice name for model
	char
	    model(namelen);


	//---------------------------------------------------------------
	//	navigation information
	//---------------------------------------------------------------
 	
     float
         staticTopo(y, x) ;
             staticTopo:units = "meters";
             staticTopo:long_name = "Topography";
             staticTopo:_FillValue = -99999.f;
     float
         staticCoriolis(y, x) ;
             staticCoriolis:units = "/second";
             staticCoriolis:long_name = "Coriolis parameter";
             staticCoriolis:_FillValue = -99999.f;
     float
         staticSpacing(y, x) ;
             staticSpacing:units = "meters";
             staticSpacing:long_name = "Grid spacing";
             staticSpacing:_FillValue = -99999.f;

// global attributes:
     :cdlDate = "20001009";
     :depictorName = "cwblaps" ;
     :projIndex = 3 ;
     :projName = "LAMBERT_CONFORMAL";
     :centralLat = 10.f ;
     :centralLon = 120.f ;
     :rotation = 40.f ;
     :xMin = -0.025650f ;
     :xMax = 0.36983f ;
     :yMax = -0.795383f ;
     :yMin = -0.873200f ;
     :lat00 = 17.8164f ;
     :lon00 = 116.065f ;
     :latNxNy = 29.18094f ;
     :lonNxNy = 126.2259f ;
     :dxKm = 5.000f ;
     :dyKm = 5.000f ;
     :latDxDy = 23.5f ;
     :lonDxDy = 121.15f ;

    data:
	origin 		= "NOAA/ERL Forecast Systems Laboratory, Boulder CO";
	model 		= "Local Analysis and Prediction System model";

	// Forecast times(hrs) are: 0(Analysis)
	valtimeMINUSreftime = 0;

        ghLevels	= "MB 1100   ",
			  "MB 1050   ",
			  "MB 1000   ",
                          "MB 950    ",
                          "MB 900    ",
                          "MB 850    ",
                          "MB 800    ",
                          "MB 750    ",
                          "MB 700    ",
                          "MB 650    ",
                          "MB 600    ",
                          "MB 550    ",
                          "MB 500    ",
                          "MB 450    ",
                          "MB 400    ",
                          "MB 350    ",
                          "MB 300    ",
                          "MB 250    ",
                          "MB 200    ",
                          "MB 150    ",
                          "MB 100    ";
        rhLevels	= "SFC       ",
			  "MB 1100   ",
			  "MB 1050   ",
			  "MB 1000   ",
                          "MB 950    ",
                          "MB 900    ",
                          "MB 850    ",
                          "MB 800    ",
                          "MB 750    ",
                          "MB 700    ",
                          "MB 650    ",
                          "MB 600    ",
                          "MB 550    ",
                          "MB 500    ",
                          "MB 450    ",
                          "MB 400    ",
                          "MB 350    ",
                          "MB 300    ",
                          "MB 250    ",
                          "MB 200    ",
                          "MB 150    ",
                          "MB 100    ";
        tLevels		= "SFC       ",
     			  "MB 1100   ",
			  "MB 1050   ",
			  "MB 1000   ",
                          "MB 950    ",
                          "MB 900    ",
                          "MB 850    ",
                          "MB 800    ",
                          "MB 750    ",
                          "MB 700    ",
                          "MB 650    ",
                          "MB 600    ",
                          "MB 550    ",
                          "MB 500    ",
                          "MB 450    ",
                          "MB 400    ",
                          "MB 350    ",
                          "MB 300    ",
                          "MB 250    ",
                          "MB 200    ",
                          "MB 150    ",
                          "MB 100    ";
        uwLevels	= "SFC       ",
			  "MB 1100   ",
			  "MB 1050   ",
			  "MB 1000   ",
                          "MB 950    ",
                          "MB 900    ",
                          "MB 850    ",
                          "MB 800    ",
                          "MB 750    ",
                          "MB 700    ",
                          "MB 650    ",
                          "MB 600    ",
                          "MB 550    ",
                          "MB 500    ",
                          "MB 450    ",
                          "MB 400    ",
                          "MB 350    ",
                          "MB 300    ",
                          "MB 250    ",
                          "MB 200    ",
                          "MB 150    ",
                          "MB 100    ";
        vwLevels	= "SFC       ",
			  "MB 1100   ",
			  "MB 1050   ",
			  "MB 1000   ",
                          "MB 950    ",
                          "MB 900    ",
                          "MB 850    ",
                          "MB 800    ",
                          "MB 750    ",
                          "MB 700    ",
                          "MB 650    ",
                          "MB 600    ",
                          "MB 550    ",
                          "MB 500    ",
                          "MB 450    ",
                          "MB 400    ",
                          "MB 350    ",
                          "MB 300    ",
                          "MB 250    ",
                          "MB 200    ",
                          "MB 150    ",
                          "MB 100    ";
       pvvLevels	= "SFC       ",
			  "MB 1100   ",
			  "MB 1050   ",
			  "MB 1000   ",
                          "MB 950    ",
                          "MB 900    ",
                          "MB 850    ",
                          "MB 800    ",
                          "MB 750    ",
                          "MB 700    ",
                          "MB 650    ",
                          "MB 600    ",
                          "MB 550    ",
                          "MB 500    ",
                          "MB 450    ",
                          "MB 400    ",
                          "MB 350    ",
                          "MB 300    ",
                          "MB 250    ",
                          "MB 200    ",
                          "MB 150    ",
                          "MB 100    ";
        shLevels	= "MB 1100   ",
			  "MB 1050   ",
			  "MB 1000   ",
                          "MB 950    ",
                          "MB 900    ",
                          "MB 850    ",
                          "MB 800    ",
                          "MB 750    ",
                          "MB 700    ",
                          "MB 650    ",
                          "MB 600    ",
                          "MB 550    ",
                          "MB 500    ",
                          "MB 450    ",
                          "MB 400    ",
                          "MB 350    ",
                          "MB 300    ",
                          "MB 250    ",
                          "MB 200    ",
                          "MB 150    ",
                          "MB 100    ";
        rrLevels	= "MB 1100   ",
			  "MB 1050   ",
			  "MB 1000   ",
                          "MB 950    ",
                          "MB 900    ",
                          "MB 850    ",
                          "MB 800    ",
                          "MB 750    ",
                          "MB 700    ",
                          "MB 650    ",
                          "MB 600    ",
                          "MB 550    ",
                          "MB 500    ",
                          "MB 450    ",
                          "MB 400    ",
                          "MB 350    ",
                          "MB 300    ",
                          "MB 250    ",
                          "MB 200    ",
                          "MB 150    ",
                          "MB 100    ";
        ptypLevels	= "MB 1100   ",
			  "MB 1050   ",
			  "MB 1000   ",
                          "MB 950    ",
                          "MB 900    ",
                          "MB 850    ",
                          "MB 800    ",
                          "MB 750    ",
                          "MB 700    ",
                          "MB 650    ",
                          "MB 600    ",
                          "MB 550    ",
                          "MB 500    ",
                          "MB 450    ",
                          "MB 400    ",
                          "MB 350    ",
                          "MB 300    ",
                          "MB 250    ",
                          "MB 200    ",
                          "MB 150    ",
                          "MB 100    ";
        ctypLevels	= "MB 1100   ",
			  "MB 1050   ",
			  "MB 1000   ",
                          "MB 950    ",
                          "MB 900    ",
                          "MB 850    ",
                          "MB 800    ",
                          "MB 750    ",
                          "MB 700    ",
                          "MB 650    ",
                          "MB 600    ",
                          "MB 550    ",
                          "MB 500    ",
                          "MB 450    ",
                          "MB 400    ",
                          "MB 350    ",
                          "MB 300    ",
                          "MB 250    ",
                          "MB 200    ",
                          "MB 150    ",
                          "MB 100    ";
        ccpcLevels	= "MB 1100   ",
			  "MB 1050   ",
			  "MB 1000   ",
                          "MB 950    ",
                          "MB 900    ",
                          "MB 850    ",
                          "MB 800    ",
                          "MB 750    ",
                          "MB 700    ",
                          "MB 650    ",
                          "MB 600    ",
                          "MB 550    ",
                          "MB 500    ",
                          "MB 450    ",
                          "MB 400    ",
                          "MB 350    ",
                          "MB 300    ",
                          "MB 250    ",
                          "MB 200    ",
                          "MB 150    ",
                          "MB 100    ";
        cwLevels	= "MB 1100   ",
			  "MB 1050   ",
			  "MB 1000   ",
                          "MB 950    ",
                          "MB 900    ",
                          "MB 850    ",
                          "MB 800    ",
                          "MB 750    ",
                          "MB 700    ",
                          "MB 650    ",
                          "MB 600    ",
                          "MB 550    ",
                          "MB 500    ",
                          "MB 450    ",
                          "MB 400    ",
                          "MB 350    ",
                          "MB 300    ",
                          "MB 250    ",
                          "MB 200    ",
                          "MB 150    ",
                          "MB 100    ";
        ciceLevels	= "MB 1100   ",
			  "MB 1050   ",
			  "MB 1000   ",
                          "MB 950    ",
                          "MB 900    ",
                          "MB 850    ",
                          "MB 800    ",
                          "MB 750    ",
                          "MB 700    ",
                          "MB 650    ",
                          "MB 600    ",
                          "MB 550    ",
                          "MB 500    ",
                          "MB 450    ",
                          "MB 400    ",
                          "MB 350    ",
                          "MB 300    ",
                          "MB 250    ",
                          "MB 200    ",
                          "MB 150    ",
                          "MB 100    ";
        hycLevels	= "MB 1100   ",
			  "MB 1050   ",
			  "MB 1000   ",
                          "MB 950    ",
                          "MB 900    ",
                          "MB 850    ",
                          "MB 800    ",
                          "MB 750    ",
                          "MB 700    ",
                          "MB 650    ",
                          "MB 600    ",
                          "MB 550    ",
                          "MB 500    ",
                          "MB 450    ",
                          "MB 400    ",
                          "MB 350    ",
                          "MB 300    ",
                          "MB 250    ",
                          "MB 200    ",
                          "MB 150    ",
                          "MB 100    ";
	pLevels		= "SFC       ",
			  "FH 1500   ";
	mslpLevels	= "SFC       ";
	dptLevels	= "SFC       ";
	potLevels	= "SFC       ";
	ccLevels	= "SFC       ",
			  "MSL       ";
	tadvLevels	= "SFC       ";
	eptLevels	= "SFC       ";
	ilwLevels	= "SFC       ";
	mconLevels	= "SFC       ";
	ptaLevels	= "SFC       ";
	sliLevels	= "SFC       ";
	hidxLevels	= "SFC       ";
	cssiLevels	= "SFC       ";
	pbeLevels	= "SFC       ";
	nbeLevels	= "SFC       ";
	visLevels	= "SFC       ";
	ccovLevels	= "SFC       ";
	cbLevels	= "SFC       ";
	ctopLevels	= "SFC       ";
	mretLevels	= "SFC       ";
	llrLevels	= "SFC       ";
	heliLevels	= "SFC       ";
	tpwLevels	= "SFC       ";
	s1hrLevels	= "SFC       ";
	stotLevels	= "SFC       ";
	pcLevels	= "SFC       ";
	stpaLevels	= "SFC       ";
	sptLevels	= "SFC       ";
	pttLevels	= "SFC       ";
	fdLevels	= "SFC       ";
	scpLevels	= "SFC       ";
	smcLevels	= "BLS  1    ",
			  "BLS  2    ",
		 	  "BLS  3    ";
}


