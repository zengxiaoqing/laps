netcdf lvd {

    dimensions:
        record = unlimited,
        z = 1,
	x = 125,
	y = 105,
        nav = 1,
        namelen = 132;
		
    variables:
        //	satellite IR channel 4 b-temp: warmest pixl

	float                                  
            s8w(record,z,y,x);
            s8w:navigation_dim = "nav";
            s8w:record = "valtime, reftime";
            s8w:_FillValue = 1.e+37f;
            s8w:long_name="IR channel 4 (11.2u) b-temp: warmest pixel";
            s8w:units="degrees Kelvin";
            s8w:valid_range= 0.f, 400.f;
            s8w:LAPS_var="S8W";
            s8w:lvl_coord=" ";
            s8w:LAPS_units="K";
                	        
        //	satellite IR channel 4 b-temp: coldest pixl

	float                                  
            s8c(record,z,y,x);
            s8c:navigation_dim = "nav";
            s8c:record = "valtime, reftime";
            s8c:_FillValue = 1.e+37f;
            s8c:long_name="IR channel 4 (11.2u) b-temp: coldest pixel";
            s8c:units="degrees Kelvin";
            s8c:valid_range= 0.f, 400.f;
            s8c:LAPS_var="S8C";
            s8c:lvl_coord=" ";
            s8c:LAPS_units="K";
                	        
        //	satellite vis counts - raw 

	float                                  
            svs(record,z,y,x);
            svs:navigation_dim = "nav";
            svs:record = "valtime, reftime";
            svs:_FillValue = 1.e+37f;
            svs:long_name="visible satellite counts - raw";
            svs:units="counts";
            svs:valid_range= 0, 3;
            svs:LAPS_var="SVS";
            svs:lvl_coord="   ";
            svs:LAPS_units="COUNTS";
                	        
        //	 satellite vis counts - normalized

	float                                  
            svn(record,z,y,x);
            svn:navigation_dim = "nav";
            svn:record = "valtime, reftime";
            svn:_FillValue = 1.e+37f;
            svn:long_name="visible satellite counts - normalized";
            svn:units="counts";
            svn:valid_range= 0, 255;
            svn:LAPS_var="SVN";
            svn:lvl_coord=" ";
            svn:LAPS_units="COUNTS";
                	        
        //	laps-albedo

	float                                  
            alb(record,z,y,x);
            alb:navigation_dim = "nav";
            alb:record = "valtime, reftime";
            alb:_FillValue = 1.e+37f;
            alb:long_name="laps derived albedo";
            alb:units="none";
            alb:valid_range= -1.f, 1.f;
            alb:LAPS_var="ALB";
            alb:lvl_coord=" ";
            alb:LAPS_units=" ";
                	        
        //	satellite IR channel 2 b-temp: averaged

	float                                  
            s3a(record,z,y,x);
            s3a:navigation_dim = "nav";
            s3a:record = "valtime, reftime";
            s3a:_FillValue = 1.e+37f;
            s3a:long_name="IR channel 2 (3.9u) b-temp: averaged";
            s3a:units="degrees Kelvin";
            s3a:valid_range= 0.f, 400.f;
            s3a:LAPS_var="S3A";
            s3a:lvl_coord=" ";
            s3a:LAPS_units="K";
                	        
        //	satellite IR channel 2 b-temp: filtered

	float                                  
            s3c(record,z,y,x);
            s3c:navigation_dim = "nav";
            s3c:record = "valtime, reftime";
            s3c:_FillValue = 1.e+37f;
            s3c:long_name="IR channel 2 (3.9u) b-temp: filtered";
            s3c:units="degrees Kelvin";
            s3c:valid_range= 0.f, 400.f;
            s3c:LAPS_var="S3C";
            s3c:lvl_coord=" ";
            s3c:LAPS_units="K";

        //	satellite IR channel 3 b-temp: averaged	

	float                                  
            s4a(record,z,y,x);
            s4a:navigation_dim = "nav";
            s4a:record = "valtime, reftime";
            s4a:_FillValue = 1.e+37f;
            s4a:long_name="IR channel 3 (6.7u) b-temp: averaged";
            s4a:units="degrees Kelvin";
            s4a:valid_range= 0.f, 400.f;
            s4a:LAPS_var="S4A";
            s4a:lvl_coord=" ";
            s4a:LAPS_units="K";

        //	satellite IR channel 3 b-temp: filtered

	float                                  
            s4c(record,z,y,x);
            s4c:navigation_dim = "nav";
            s4c:record = "valtime, reftime";
            s4c:_FillValue = 1.e+37f;
            s4c:long_name="IR channel 3 (6.7u) b-temp: filtered";
            s4c:units="degrees Kelvin";
            s4c:valid_range= 0.f, 400.f;
            s4c:LAPS_var="S4C";
            s4c:lvl_coord=" ";
            s4c:LAPS_units="K";

        //	satellite IR unused

	float                                  
            s5a(record,z,y,x);
            s5a:navigation_dim = "nav";
            s5a:record = "valtime, reftime";
            s5a:_FillValue = 1.e+37f;
            s5a:long_name="unused";
            s5a:units="degrees Kelvin";
            s5a:valid_range= 0.f, 400.f;
            s5a:LAPS_var="S5A";
            s5a:lvl_coord=" ";
            s5a:LAPS_units="K";

        //	satellite IR unused

	float                                  
            s5c(record,z,y,x);
            s5c:navigation_dim = "nav";
            s5c:record = "valtime, reftime";
            s5c:_FillValue = 1.e+37f;
            s5c:long_name="unused";
            s5c:units="degrees Kelvin";
            s5c:valid_range= 0.f, 400.f;
            s5c:LAPS_var="S5C";
            s5c:lvl_coord=" ";
            s5c:LAPS_units="K";

        //	 satellite IR channel 4 b-temp: averaged

	float                                  
            s8a(record,z,y,x);
            s8a:navigation_dim = "nav";
            s8a:record = "valtime, reftime";
            s8a:_FillValue = 1.e+37f;
            s8a:long_name="IR channel 4 (11.2u) b-temp: averaged";
            s8a:units="degrees Kelvin";
            s8a:valid_range= 0.f, 400.f;
            s8a:LAPS_var="S8A";
            s8a:lvl_coord=" ";
            s8a:LAPS_units="K";

        //	satellite IR channel 5 b-temp: averaged

	float                                  
            sca(record,z,y,x);
            sca:navigation_dim = "nav";
            sca:record = "valtime, reftime";
            sca:_FillValue = 1.e+37f;
            sca:long_name="IR channel 5 (12.0u) b-temp: averaged";
            sca:units="degrees Kelvin";
            sca:valid_range= 0.f, 400.f;
            sca:LAPS_var="SCA";
            sca:lvl_coord=" ";
            sca:LAPS_units="K";

        //	satellite IR channel 5 b-temp: filtered

	float                                  
            scc(record,z,y,x);
            scc:navigation_dim = "nav";
            scc:record = "valtime, reftime";
            scc:_FillValue = 1.e+37f;
            scc:long_name="IR channel 5 (12.0u) b-temp: filtered";
            scc:units="degrees Kelvin";
            scc:valid_range= 0.f, 400.f;
            scc:LAPS_var="SCC";
            scc:lvl_coord=" ";
            scc:LAPS_units="K";

        //	LAPS variables

        long
            imax,
            jmax,
            kmax,
            kdim;

        char
            s8w_comment(record,z,namelen),
            s8c_comment(record,z,namelen),
            svs_comment(record,z,namelen),
            svn_comment(record,z,namelen),
            alb_comment(record,z,namelen),
            s3a_comment(record,z,namelen),
            s3c_comment(record,z,namelen),
            s4a_comment(record,z,namelen),
            s4c_comment(record,z,namelen),
            s5a_comment(record,z,namelen),
            s5c_comment(record,z,namelen),
            s8a_comment(record,z,namelen),
            sca_comment(record,z,namelen),
            scc_comment(record,z,namelen),
            asctime(record,namelen);

			
        //	inventory variables

        short
            s8w_fcinv(record, z);
            s8w_fcinv:_FillValue= 0s;
              	
        short
            s8c_fcinv(record, z);
            s8c_fcinv:_FillValue= 0s;
              	
        short
            svs_fcinv(record, z);
            svs_fcinv:_FillValue= 0s;
              	
        short
            svn_fcinv(record, z);
            svn_fcinv:_FillValue= 0s;
              	
        short
            alb_fcinv(record, z);
            alb_fcinv:_FillValue= 0s;
              	
        short
            s3a_fcinv(record, z);
            s3a_fcinv:_FillValue= 0s;
              	
        short
            s3c_fcinv(record, z);
            s3c_fcinv:_FillValue= 0s;
              	
        short
            s4a_fcinv(record, z);
            s4a_fcinv:_FillValue= 0s;
              	
        short
            s4c_fcinv(record, z);
            s4c_fcinv:_FillValue= 0s;
              	
        short
            s5a_fcinv(record, z);
            s5a_fcinv:_FillValue= 0s;
              	
        short
            s5c_fcinv(record, z);
            s5c_fcinv:_FillValue= 0s;
              	
        short
            s8a_fcinv(record, z);
            s8a_fcinv:_FillValue= 0s;
              	
        short
            sca_fcinv(record, z);
            sca_fcinv:_FillValue= 0s;
              	
        short
            scc_fcinv(record, z);
            scc_fcinv:_FillValue= 0s;
              	
        //	list of grid levels

        float 
            level(z);
            level:long_name="level of data";
	    level:units = "hectopascals";
                    	
        //      validtime of the grid 

        double
            valtime(record);
            valtime:long_name = "valid time";
            valtime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      reference time of the process

        double
            reftime(record);
            reftime:long_name = "reference time";
            reftime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      nice name for originating center

        char
            origin_name(namelen);

        //      nice name for process

        char
            process_name(namelen);

        //      nice name for grid description instance
        char
            grid_name(namelen);

        //      basic assumption about earth shape
        char
            earth_shape(namelen);

        // navigation variables using 
        // WMO FM 92-VIII Ext.GRIB specification names
  
        char    grid_type(nav, namelen);
                grid_type:long_name = "GRIB-1 grid type";
  
        char    x_dim(nav, namelen);
                x_dim:long_name = "longitude dimension";
  
        char    y_dim(nav, namelen);
                y_dim:long_name = "latitude dimension";
  
        short   Nx(nav);
                Nx:long_name = "number of x points";
  
        short   Ny(nav);
                Ny:long_name =  "number of y points";
  
        float   La1(nav);
                La1:long_name = "first latitude";
                La1:units = "degrees_north";
  
        float   Lo1(nav);
                Lo1:long_name = "first longitude";
                Lo1:units = "degrees_east" ;
    
        float   LoV(nav);
                LoV:long_name = "orientation of grid" ;
                LoV:units = "degrees_east";
  
        float   Latin1(nav);
                Latin1:long_name = "orientation of grid" ;
                Latin1:units = "degrees_north";

        float   Latin2(nav);
                Latin2:long_name = "orientation of grid" ;
                Latin2:units = "degrees_north";

        float   Dx(nav);
                Dx:long_name = "x grid increment";
                Dx:units = "meters";
  
        float   Dy(nav);
                Dy:long_name = "y grid increment";
                Dy:units = "meters";
  
        // end of navigation variables

        :Conventions = "NUWG";
        :history = "created by LAPS Branch of FSL";
        :record = "valtime, reftime";
        :title = "LAPS lvd file - satellite data";
        :version = 3;

    data:

        earth_shape     = "spherical radius";
        grid_name       = "LAPS lvd file - satellite data";
        process_name    = "LAPS - Local Analysis and Prediction System";
        x_dim           = "x";
        y_dim           = "y";
}                       
