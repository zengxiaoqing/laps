netcdf lcb {

    dimensions:
        record = unlimited,
        z = 1,
	x = 125,
	y = 105,
        nav = 1,
        namelen = 132;
		
    variables:
        //	cloud base

	float                                  
            lcb(record,z,y,x);
            lcb:navigation_dim = "nav";
            lcb:record = "valtime, reftime";
            lcb:_FillValue = 1.e+37f;
            lcb:long_name="LAPS cloud base";
            lcb:units="meters";
            lcb:valid_range= -200.f, 200.f;
            lcb:LAPS_var="LCB";
            lcb:lvl_coord="MSL";
	    lcb:LAPS_units="M";
                	        
        //	cloud top

	float                                  
            lct(record,z,y,x);
            lct:navigation_dim = "nav";
            lct:record = "valtime, reftime";
            lct:_FillValue = 1.e+37f;
            lct:long_name="LAPS cloud top";
            lct:units="meters";
            lct:valid_range= -200.f, 200.f;
            lct:LAPS_var="LCT";
            lct:lvl_coord="MSL";
	    lct:LAPS_units="M";
                	        
        //	cloud ceiling 
        float 
            cce(record,z,y,x) ;
            cce:navigation_dim = "nav";
            cce:record = "valtime, reftime";
            cce:_FillValue = 1.e+37f;
            cce:long_name="LAPS cloud ceiling" ;
            cce:units = "meters" ;
            cce:valid_range = 0.f, 40000.f ;
            cce:LAPS_var = "CCE" ;
            cce:lvl_coord = "AGL" ;
            cce:LAPS_units = "M" ;
                	        
        //	cloud parallax 
        float 
            plx(record,z,y,x) ;
            plx:navigation_dim = "nav";
            plx:record = "valtime, reftime";
            plx:_FillValue = 1.e+37f;
            plx:long_name="cloud parallax" ;
            plx:units = "meters" ;
            plx:valid_range = 0.f, 40000.f ;
            plx:LAPS_var = "PLX" ;
            plx:lvl_coord = " " ;
            plx:LAPS_units = "M" ;


        //	LAPS variables

        long
            imax,
            jmax,
            kmax,
            kdim;

        char
            lcb_comment(record,z,namelen),
            lct_comment(record,z,namelen),
            cce_comment(record,z,namelen),
            plx_comment(record,z,namelen),
            asctime(record,namelen);

			
        //	inventory variables

        short
            lcb_fcinv(record, z);
            lcb_fcinv:_FillValue= 0s;
              	
        short
            lct_fcinv(record, z);
            lct_fcinv:_FillValue= 0s;
              	
        short
            cce_fcinv(record, z);
            cce_fcinv:_FillValue= 0s;
              	
        short
            plx_fcinv(record, z);
            plx_fcinv:_FillValue= 0s;
              	
        //	list of grid levels

        float 
            level(z);
            level:long_name="level of data";
	    level:units = "hectopascals";
                    	
        //      validtime of the grid 

        double
            valtime(record);
            valtime:long_name = "valid time";
            valtime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      reference time of the process

        double
            reftime(record);
            reftime:long_name = "reference time";
            reftime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      nice name for originating center

        char
            origin_name(namelen);

        //      nice name for process

        char
            process_name(namelen);

        //      nice name for grid description instance
        char
            grid_name(namelen);

        //      basic assumption about earth shape
        char
            earth_shape(namelen);

        // navigation variables using 
        // WMO FM 92-VIII Ext.GRIB specification names
  
        char    grid_type(nav, namelen);
                grid_type:long_name = "GRIB-1 grid type";
  
        char    x_dim(nav, namelen);
                x_dim:long_name = "longitude dimension";
  
        char    y_dim(nav, namelen);
                y_dim:long_name = "latitude dimension";
  
        short   Nx(nav);
                Nx:long_name = "number of x points";
  
        short   Ny(nav);
                Ny:long_name =  "number of y points";
  
        float   La1(nav);
                La1:long_name = "first latitude";
                La1:units = "degrees_north";
  
        float   Lo1(nav);
                Lo1:long_name = "first longitude";
                Lo1:units = "degrees_east" ;
    
        float   LoV(nav);
                LoV:long_name = "orientation of grid" ;
                LoV:units = "degrees_east";
  
        float   Latin1(nav);
                Latin1:long_name = "orientation of grid" ;
                Latin1:units = "degrees_north";

        float   Latin2(nav);
                Latin2:long_name = "orientation of grid" ;
                Latin2:units = "degrees_north";

        float   Dx(nav);
                Dx:long_name = "x grid increment";
                Dx:units = "meters";
  
        float   Dy(nav);
                Dy:long_name = "y grid increment";
                Dy:units = "meters";
  
        // end of navigation variables

        :Conventions = "NUWG";
        :history = "created by LAPS Branch of FSL";
        :record = "valtime, reftime";
        :title = "LAPS lcb file - LAPS cloud base and top";
        :version = 3;

    data:

        earth_shape     = "spherical radius";
        grid_name       = "LAPS lcb file - LAPS cloud base and top";
        process_name    = "LAPS - Local Analysis and Prediction System";
        x_dim           = "x";
        y_dim           = "y";
}                       
