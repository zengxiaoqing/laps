netcdf ln3 {

    dimensions:
        record = unlimited,
        z = 1,
	x = 125,
	y = 105,
        nav = 1,
        namelen = 132;
		
    variables:
        //	3D radar - low level layer composite reflectivity

	float                                  
            r04(record,z,y,x);
            r04:navigation_dim = "nav";
            r04:record = "valtime, reftime";
            r04:_FillValue = 1.e+37f;
            r04:long_name="low level layer composite reflectivity";
            r04:units="dBZ";
            r04:valid_range= -10.f, 80.f;
            r04:LAPS_var="R04";
            r04:lvl_coord="    ";
	    r04:LAPS_units="DBZ       ";
                	        
        //	3D radar - mid level layer composite reflectivity

	float                                  
            r48(record,z,y,x);
            r48:navigation_dim = "nav";
            r48:record = "valtime, reftime";
            r48:_FillValue = 1.e+37f;
            r48:long_name="mid level layer composite reflectivity";
            r48:units="dBZ";
            r48:valid_range= -10.f, 80.f;
            r48:LAPS_var="R48";
            r48:lvl_coord="    ";
	    r48:LAPS_units="DBZ       ";
               	        
        //	3D radar - high level layer composite reflectivity

	float                                  
            r8c(record,z,y,x);
            r8c:navigation_dim = "nav";
            r8c:record = "valtime, reftime";
            r8c:_FillValue = 1.e+37f;
            r8c:long_name="high level layer composite reflectivity";
            r8c:units="dBZ";
            r8c:valid_range= -10.f, 80.f;
            r8c:LAPS_var="R8C";
            r8c:lvl_coord="    ";
	    r8c:LAPS_units="DBZ       ";
                	        
        //	3D radar - echo tops height

	float                                  
            et(record,z,y,x);
            et:navigation_dim = "nav";
            et:record = "valtime, reftime";
            et:_FillValue = 1.e+37f;
            et:long_name="echo tops height";
            et:units="meters";
            et:valid_range= 0.f, 30000.f;
            et:LAPS_var="ET ";
            et:lvl_coord="MSL ";
	    et:LAPS_units="M         ";
                	        
        //	3D radar - composite reflectivity

	float                                  
            rco(record,z,y,x);
            rco:navigation_dim = "nav";
            rco:record = "valtime, reftime";
            rco:_FillValue = 1.e+37f;
            rco:long_name="composite reflectivity";
            rco:units="dBZ";
            rco:valid_range= -10.f, 80.f;
            rco:LAPS_var="RCO";
            rco:lvl_coord="    ";
	    rco:LAPS_units="DBZ       ";
                	        
        //	3D radar - radar vertically integrated liquid

	float                                  
            vil(record,z,y,x);
            vil:navigation_dim = "nav";
            vil:record = "valtime, reftime";
            vil:_FillValue = 1.e+37f;
            vil:long_name="radar vertically integrated liquid";
            vil:units="grams/meter**2";
            vil:valid_range= 0.f, 0.1f;
            vil:LAPS_var="VIL";
            vil:lvl_coord="    ";
	    vil:LAPS_units="G/M**2    ";
                	        
        //	LAPS variables

        long
            imax,
            jmax,
            kmax,
            kdim;

        char
            r04_comment(record,z,namelen),
            r48_comment(record,z,namelen),
            r8c_comment(record,z,namelen),
            et_comment(record,z,namelen),
            rco_comment(record,z,namelen),
            vil_comment(record,z,namelen),
            asctime(record,namelen);

			
        //	inventory variables

        short
            r04_fcinv(record, z);
            r04_fcinv:_FillValue= 0s;
              	
        short
            r48_fcinv(record, z);
            r48_fcinv:_FillValue= 0s;
              	
        short
            r8c_fcinv(record, z);
            r8c_fcinv:_FillValue= 0s;
              	
        short
            et_fcinv(record, z);
            et_fcinv:_FillValue= 0s;
              	
        short
            rco_fcinv(record, z);
            rco_fcinv:_FillValue= 0s;
              	
        short
            vil_fcinv(record, z);
            vil_fcinv:_FillValue= 0s;
              	
        //	list of grid levels

        float 
            level(z);
            level:long_name="level of data";
	    level:units = "hectopascals";
                    	
        //      validtime of the grid 

        double
            valtime(record);
            valtime:long_name = "valid time";
            valtime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      reference time of the process

        double
            reftime(record);
            reftime:long_name = "reference time";
            reftime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      nice name for originating center

        char
            origin_name(namelen);

        //      nice name for process

        char
            process_name(namelen);

        //      nice name for grid description instance
        char
            grid_name(namelen);

        //      basic assumption about earth shape
        char
            earth_shape(namelen);

        // navigation variables using 
        // WMO FM 92-VIII Ext.GRIB specification names
  
        char    grid_type(nav, namelen);
                grid_type:long_name = "GRIB-1 grid type";
  
        char    x_dim(nav, namelen);
                x_dim:long_name = "longitude dimension";
  
        char    y_dim(nav, namelen);
                y_dim:long_name = "latitude dimension";
  
        short   Nx(nav);
                Nx:long_name = "number of x points";
  
        short   Ny(nav);
                Ny:long_name =  "number of y points";
  
        float   La1(nav);
                La1:long_name = "first latitude";
                La1:units = "degrees_north";
  
        float   Lo1(nav);
                Lo1:long_name = "first longitude";
                Lo1:units = "degrees_east" ;
    
        float   LoV(nav);
                LoV:long_name = "orientation of grid" ;
                LoV:units = "degrees_east";
  
        float   Latin1(nav);
                Latin1:long_name = "orientation of grid" ;
                Latin1:units = "degrees_north";

        float   Latin2(nav);
                Latin2:long_name = "orientation of grid" ;
                Latin2:units = "degrees_north";

        float   Dx(nav);
                Dx:long_name = "x grid increment";
                Dx:units = "kilometers";
  
        float   Dy(nav);
                Dy:long_name = "y grid increment";
                Dy:units = "kilometers";
  
        // end of navigation variables

        :Conventions = "NUWG";
        :history = "created by LAPS Branch of FSL";
        :record = "valtime, reftime";
        :title = "LAPS ln3 file - 3D radar";
        :version = 3;

    data:

        earth_shape     = "spherical radius";
        grid_name       = "LAPS ln3 file - 3D radar";
        process_name    = "LAPS - Local Analysis and Prediction System";
        x_dim           = "x";
        y_dim           = "y";
}                       
