netcdf lil {

    dimensions:
        record = unlimited,
        z = 1,
	x = 125,
	y = 105,
        nav = 1,
        namelen = 132;
		
    variables:
        //	integrated cloud liquid

	float                                  
            lil(record,z,y,x);
            lil:navigation_dim = "nav";
            lil:record = "valtime, reftime";
            lil:_FillValue = 1.e+37f;
            lil:long_name="integrated cloud liquid";
            lil:units="meters";
            lil:valid_range= 0.f, 100.f;
            lil:LAPS_var="LIL";
            lil:lvl_coord="MSL";
	    lil:LAPS_units="M";

        //	integrated cloud ice               

	float                                  
            lic(record,z,y,x);
            lic:navigation_dim = "nav";
            lic:record = "valtime, reftime";
            lic:_FillValue = 1.e+37f;
            lic:long_name="integrated cloud ice";
            lic:units="meters";
            lic:valid_range= 0.f, 100.f;
            lic:LAPS_var="LIC";
            lic:lvl_coord="MSL";
	    lic:LAPS_units="M";

        //	cloud optical depth

	float                                  
            cod(record,z,y,x);
            cod:navigation_dim = "nav";
            cod:record = "valtime, reftime";
            cod:_FillValue = 1.e+37f;
            cod:long_name="cloud optical depth";
            cod:units="none";
            cod:valid_range= 0.f, 1000.f;
            cod:LAPS_var="COD";
            cod:lvl_coord="MSL";
	    cod:LAPS_units="NONE";

        //      cloud albedo

        float
            cla(record,z,y,x);
            cla:_FillValue = 1.e+37f;
            cla:long_name="Cloud Albedo";
            cla:units="none";
            cla:valid_range= 0.f, 1.f;
            cla:LAPS_var="CLA";
            cla:lvl_coord="MSL";
            cla:LAPS_units="none";

        //	LAPS variables

        long
            imax,
            jmax,
            kmax,
            kdim;

        char
            lil_comment(record,z,namelen),
            lic_comment(record,z,namelen),
            cod_comment(record,z,namelen),
            cla_comment(record,z,namelen),
            asctime(record,namelen);

			
        //	inventory variables

        short
            lil_fcinv(record, z);
            lil_fcinv:_FillValue= 0s;

        short
            lic_fcinv(record, z);
            lic_fcinv:_FillValue= 0s;

        short
            cod_fcinv(record, z);
            cod_fcinv:_FillValue= 0s;

        short
            cla_fcinv(record, z);
            cla_fcinv:_FillValue= 0s;
              	
        //	list of grid levels

        float 
            level(z);
            level:long_name="level of data";
	    level:units = "hectopascals";
                    	
        //      validtime of the grid 

        double
            valtime(record);
            valtime:long_name = "valid time";
            valtime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      reference time of the process

        double
            reftime(record);
            reftime:long_name = "reference time";
            reftime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      nice name for originating center

        char
            origin_name(namelen);

        //      nice name for process

        char
            process_name(namelen);

        //      nice name for grid description instance
        char
            grid_name(namelen);

        //      basic assumption about earth shape
        char
            earth_shape(namelen);

        // navigation variables using 
        // WMO FM 92-VIII Ext.GRIB specification names
  
        char    grid_type(nav, namelen);
                grid_type:long_name = "GRIB-1 grid type";
  
        char    x_dim(nav, namelen);
                x_dim:long_name = "longitude dimension";
  
        char    y_dim(nav, namelen);
                y_dim:long_name = "latitude dimension";
  
        short   Nx(nav);
                Nx:long_name = "number of x points";
  
        short   Ny(nav);
                Ny:long_name =  "number of y points";
  
        float   La1(nav);
                La1:long_name = "first latitude";
                La1:units = "degrees_north";
  
        float   Lo1(nav);
                Lo1:long_name = "first longitude";
                Lo1:units = "degrees_east" ;
    
        float   LoV(nav);
                LoV:long_name = "orientation of grid" ;
                LoV:units = "degrees_east";
  
        float   Latin1(nav);
                Latin1:long_name = "orientation of grid" ;
                Latin1:units = "degrees_north";

        float   Latin2(nav);
                Latin2:long_name = "orientation of grid" ;
                Latin2:units = "degrees_north";

        float   Dx(nav);
                Dx:long_name = "x grid increment";
                Dx:units = "meters";
  
        float   Dy(nav);
                Dy:long_name = "y grid increment";
                Dy:units = "meters";
  
        // end of navigation variables

        :Conventions = "NUWG";
        :history = "created by LAPS Branch of FSL";
        :record = "valtime, reftime";
        :title = "LAPS lil file - integrated liquid water";
        :version = 3;

    data:

        earth_shape     = "spherical radius";
        grid_name       = "LAPS lil file - integrated liquid water";
        process_name    = "LAPS - Local Analysis and Prediction System";
        x_dim           = "x";
        y_dim           = "y";
}                       
