netcdf lcv {

    dimensions:
        record = unlimited,
        z = 1,
	x = 125,
	y = 105,
        nav = 1,
        namelen = 132;
		
    variables:
        //	LAPS cloud cover

	float                                  
            lcv(record,z,y,x);
            lcv:navigation_dim = "nav";
            lcv:record = "valtime, reftime";
            lcv:_FillValue = 1.e+37f;
            lcv:long_name="LAPS cloud cover";
            lcv:units="none";
            lcv:valid_range= 0.f, 100.f;
            lcv:LAPS_var="LCV";
            lcv:lvl_coord="MSL";
	    lcv:LAPS_units="UNDIM";
                	        
        //	Cloud analysis implied snow cover 

	float                                  
            csc(record,z,y,x);
            csc:navigation_dim = "nav";
            csc:record = "valtime, reftime";
            csc:_FillValue = 1.e+37f;
            csc:long_name="Cloud analysis implied snow cover";
            csc:units="none";
            csc:valid_range= 0.f, 1.0f;
            csc:LAPS_var="CSC";
            csc:lvl_coord="MSL";
	    csc:LAPS_units="UNDIM";
                	        
        //	Cloud analysis implied snow cover 
        float 
            cwt(record,z,y,x) ;
            cwt:navigation_dim = "nav";
            cwt:record = "valtime, reftime";
            cwt:_FillValue = 1.e+37f;
            cwt:long_name = "Clear Sky Water Temperature" ;
            cwt:units = "none" ;
            cwt:valid_range = 100.f, 366.f ;
            cwt:LAPS_var = "CWT" ;
            cwt:lvl_coord = "MSL" ;
            cwt:LAPS_units = "UNDIM" ;

        //	LAPS variables

        long
            imax,
            jmax,
            kmax,
            kdim;

        char
            lcv_comment(record,z,namelen),
            csc_comment(record,z,namelen),
            cwt_comment(record,z,namelen),
            asctime(record,namelen);

			
        //	inventory variables

        short
            lcv_fcinv(record, z);
            lcv_fcinv:_FillValue= 0s;
              	
        short
            csc_fcinv(record, z);
            csc_fcinv:_FillValue= 0s;
              	
        short
            cwt_fcinv(record, z);
            cwt_fcinv:_FillValue= 0s;
              	
        //	list of grid levels

        float 
            level(z);
            level:long_name="level of data";
	    level:units = "hectopascals";
                    	
        //      validtime of the grid 

        double
            valtime(record);
            valtime:long_name = "valid time";
            valtime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      reference time of the process

        double
            reftime(record);
            reftime:long_name = "reference time";
            reftime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      nice name for originating center

        char
            origin_name(namelen);

        //      nice name for process

        char
            process_name(namelen);

        //      nice name for grid description instance
        char
            grid_name(namelen);

        //      basic assumption about earth shape
        char
            earth_shape(namelen);

        // navigation variables using 
        // WMO FM 92-VIII Ext.GRIB specification names
  
        char    grid_type(nav, namelen);
                grid_type:long_name = "GRIB-1 grid type";
  
        char    x_dim(nav, namelen);
                x_dim:long_name = "longitude dimension";
  
        char    y_dim(nav, namelen);
                y_dim:long_name = "latitude dimension";
  
        short   Nx(nav);
                Nx:long_name = "number of x points";
  
        short   Ny(nav);
                Ny:long_name =  "number of y points";
  
        float   La1(nav);
                La1:long_name = "first latitude";
                La1:units = "degrees_north";
  
        float   Lo1(nav);
                Lo1:long_name = "first longitude";
                Lo1:units = "degrees_east" ;
    
        float   LoV(nav);
                LoV:long_name = "orientation of grid" ;
                LoV:units = "degrees_east";
  
        float   Latin1(nav);
                Latin1:long_name = "orientation of grid" ;
                Latin1:units = "degrees_north";

        float   Latin2(nav);
                Latin2:long_name = "orientation of grid" ;
                Latin2:units = "degrees_north";

        float   Dx(nav);
                Dx:long_name = "x grid increment";
                Dx:units = "kilometers";
  
        float   Dy(nav);
                Dy:long_name = "y grid increment";
                Dy:units = "kilometers";
  
        // end of navigation variables

        :Conventions = "NUWG";
        :history = "created by LAPS Branch of FSL";
        :record = "valtime, reftime";
        :title = "LAPS lcv file - LAPS cloud and snow cover";
        :version = 3;

    data:

        earth_shape     = "spherical radius";
        grid_name       = "LAPS lcv file - LAPS cloud and snow cover";
        process_name    = "LAPS - Local Analysis and Prediction System";
        x_dim           = "x";
        y_dim           = "y";
}                       
