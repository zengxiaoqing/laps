netcdf lty {

    dimensions:
        record = unlimited,
        z = 21,
	x = 125,
	y = 105,
        nav = 1,
        namelen = 132;
		
    variables:
        //	precipitation type

	float                                  
            pty(record,z,y,x);
            pty:navigation_dim = "nav";
            pty:record = "valtime, reftime";
            pty:_FillValue = 1.e+37f;
            pty:long_name="precipitation type";
            pty:units="none";
            pty:valid_range= -200.f, 200.f;
            pty:LAPS_var="PTY";
            pty:lvl_coord="HPA";
	    pty:LAPS_units="NONE";
                	        
        //	cloud type

	float                                  
            cty(record,z,y,x);
            cty:navigation_dim = "nav";
            cty:record = "valtime, reftime";
            cty:_FillValue = 1.e+37f;
            cty:long_name="cloud type";
            cty:units="none";
            cty:valid_range= -200.f, 200.f;
            cty:LAPS_var="CTY";
            cty:lvl_coord="HPA";
	    cty:LAPS_units="NONE";
                	        
        //	LAPS variables

        long
            imax,
            jmax,
            kmax,
            kdim;

        char
            pty_comment(record,z,namelen),
            cty_comment(record,z,namelen),
            asctime(record,namelen);

			
        //	inventory variables

        short
            pty_fcinv(record, z);
            pty_fcinv:_FillValue= 0s;
              	
        short
            cty_fcinv(record, z);
            cty_fcinv:_FillValue= 0s;
              	
        //	list of grid levels

        float 
            level(z);
            level:long_name="level of data";
	    level:units = "hectopascals";
                    	
        //      validtime of the grid 

        double
            valtime(record);
            valtime:long_name = "valid time";
            valtime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      reference time of the process

        double
            reftime(record);
            reftime:long_name = "reference time";
            reftime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      nice name for originating center

        char
            origin_name(namelen);

        //      nice name for process

        char
            process_name(namelen);

        //      nice name for grid description instance
        char
            grid_name(namelen);

        //      basic assumption about earth shape
        char
            earth_shape(namelen);

        // navigation variables using 
        // WMO FM 92-VIII Ext.GRIB specification names
  
        char    grid_type(nav, namelen);
                grid_type:long_name = "GRIB-1 grid type";
  
        char    x_dim(nav, namelen);
                x_dim:long_name = "longitude dimension";
  
        char    y_dim(nav, namelen);
                y_dim:long_name = "latitude dimension";
  
        short   Nx(nav);
                Nx:long_name = "number of x points";
  
        short   Ny(nav);
                Ny:long_name =  "number of y points";
  
        float   La1(nav);
                La1:long_name = "first latitude";
                La1:units = "degrees_north";
  
        float   Lo1(nav);
                Lo1:long_name = "first longitude";
                Lo1:units = "degrees_east" ;
    
        float   LoV(nav);
                LoV:long_name = "orientation of grid" ;
                LoV:units = "degrees_east";
  
        float   Latin1(nav);
                Latin1:long_name = "orientation of grid" ;
                Latin1:units = "degrees_north";

        float   Latin2(nav);
                Latin2:long_name = "orientation of grid" ;
                Latin2:units = "degrees_north";

        float   Dx(nav);
                Dx:long_name = "x grid increment";
                Dx:units = "meters";
  
        float   Dy(nav);
                Dy:long_name = "y grid increment";
                Dy:units = "meters";
  
        // end of navigation variables

        :Conventions = "NUWG";
        :history = "created by LAPS Branch of FSL";
        :record = "valtime, reftime";
        :title = "LAPS lty file - cloud and precipitation type";
        :version = 3;

    data:

        earth_shape     = "spherical radius";
        grid_name       = "LAPS lty file - cloud and precipitation type";
        process_name    = "LAPS - Local Analysis and Prediction System";
        x_dim           = "x";
        y_dim           = "y";
}                       
