netcdf fsf {

    dimensions:
        record = unlimited,
        z = 1,
	x =125,
	y = 105,
        nav = 1,
        namelen = 132;
		
    variables:

        //	LAPS Fcst sfc u wind component
        //      bigfile name = uw
	float                                  
            u(record,z,y,x);
            u:_FillValue = 1.e+37f;
            u:long_name="LAPS Fcst sfc u wind component";
            u:units="m/s";
            u:valid_range= -200.f, 200.f;
            u:LAPS_var="U";
            u:lvl_coord="AGL";
	    u:LAPS_units="M/S";
                	        
        //	LAPS Fcst sfc v wind component
        //      bigfile name = vw
	float                                  
            v(record,z,y,x);
            v:_FillValue = 1.e+37f;
            v:long_name="LAPS Fcst sfc v wind component";
            v:units="m/s";
            v:valid_range= -200.f, 200.f;
            v:LAPS_var="V";
            v:lvl_coord="AGL";
	    v:LAPS_units="M/S";
                	        
        //	LAPS Fcst sfc w wind component
        //      bigfile name = ww
	float                                  
            w(record,z,y,x);
            w:_FillValue = 1.e+37f;
            w:long_name="LAPS Fcst sfc w wind component";
            w:units="m/s";
            w:valid_range= -100.f, 100.f;
            w:LAPS_var="W";
            w:lvl_coord="AGL";
	    w:LAPS_units="M/S";
                	        
        //	LAPS Fcst sfc temperature
        //      bigfile name = t
	float                                  
            t(record,z,y,x);
            t:_FillValue = 1.e+37f;
            t:long_name="LAPS Fcst sfc temperature";
            t:units="Kelvins";
            t:valid_range= 0.f, 500.f;
            t:LAPS_var="T";
            t:lvl_coord="AGL";
	    t:LAPS_units="K";
                	        
        //	LAPS Fcst surface dewpoint
        //      bigfile name = dpt
	float                                  
            td(record,z,y,x);
            td:_FillValue = 1.e+37f;
            td:long_name="LAPS Fcst sfc dewpoint";
            td:units="Kelvins";
            td:valid_range= 0.f, 500.f;
            td:LAPS_var="TD";
            td:lvl_coord="AGL";
	    td:LAPS_units="K";

        //      LAPS Fcst relative humidity       //
        //      bigfile name = rh
        float
            rh(record,z,y,x);
            rh:_FillValue = 1.e+37f;
            rh:long_name="LAPS Fcst sfc relative humidity";
            rh:units="meters";
            rh:valid_range= 0.f, 100.f;
            rh:LAPS_var="RH";
            rh:lvl_coord="AGL";
            rh:LAPS_units="PERCENT";

        //      LAPS Fcst cloud base
        //      bigfile name = cb
        float
            lcb(record,z,y,x);
            lcb:_FillValue = 1.e+37f;
            lcb:long_name="LAPS Fcst cloud base";
            lcb:units="meters";
            lcb:valid_range= 0.f, 100000.f;
            lcb:LAPS_var="LCB";
            lcb:lvl_coord="MSL";
            lcb:LAPS_units="M";

        //      LAPS Fcst cloud top
        //      bigfile name = ctop
        float
            lct(record,z,y,x);
            lct:_FillValue = 1.e+37f;
            lct:long_name="LAPS Fcst cloud top";
            lct:units="meters";
            lct:valid_range= 0.f, 100000.f;
            lct:LAPS_var="LCT";
            lct:lvl_coord="MSL";
            lct:LAPS_units="M";

        //      LAPS Fcst MSL Pressure            //
        //      bigfile name = mslp
        float
            msl(record,z,y,x);
            msl:_FillValue = 1.e+37f;
            msl:long_name="LAPS Fcst MSL pressure";
            msl:units="pascals";
            msl:valid_range= 0.f, 100000.f;
            msl:LAPS_var="MSL";
            msl:lvl_coord="MSL";
            msl:LAPS_units="PA";

        //	LAPS Fcst 1500m pressure
        //      bigfile name = p (at level "FH  1500")
	float                                  
            p(record,z,y,x);
            p:_FillValue = 1.e+37f;
            p:long_name="LAPS Fcst 1500m pressure";
            p:units="pascals";
            p:valid_range= 0.f, 100000.f;
            p:LAPS_var="P";
            p:lvl_coord="MSL";
	    p:LAPS_units="PA";
                	        
        //      LAPS Fcst surface pressure (looks like topo)      //
        //      bigfile name = p (at level "SFC")
        float
            ps(record,z,y,x);
            ps:_FillValue = 1.e+37f;
            ps:long_name="LAPS Fcst sfc pressure";
            ps:units="pascals";
            ps:valid_range= 0.f, 100000.f;
            ps:LAPS_var="PS";
            ps:lvl_coord="AGL";
            ps:LAPS_units="PA";

        //      LAPS Fcst integrated liquid water depth         
        //      bigfile name = ilw
        float
            lil(record,z,y,x);
            lil:_FillValue = 1.e+37f;
            lil:long_name="LAPS Fcst integrated liquid water depth";
            lil:units="m";
            lil:valid_range= 0.f, 1.f;
            lil:LAPS_var="LIL";
            lil:lvl_coord="AGL";
            lil:LAPS_units="M";

        //      LAPS Fcst integrated total precip water depth        
        //      bigfile name = tpw
        float
            tpw(record,z,y,x);
            tpw:_FillValue = 1.e+37f;
            tpw:long_name="LAPS Fcst precipitable water depth";
            tpw:units="m";
            tpw:valid_range= 0.f, 1.f;
            tpw:LAPS_var="TPW";
            tpw:lvl_coord="AGL";
            tpw:LAPS_units="M";

        //      LAPS Fcst increment precip accumulation depth        
        //      bigfile name = pc
        float
            r01(record,z,y,x);
            r01:_FillValue = 1.e+37f;
            r01:long_name="LAPS Fcst increment precip accum depth";
            r01:units="m";
            r01:valid_range= 0.f, 1.f;
            r01:LAPS_var="R01";
            r01:lvl_coord="AGL";
            r01:LAPS_units="M";

        //      LAPS Fcst storm total precip accumulation depth        
        //      bigfile name = stpa
        float
            rto(record,z,y,x);
            rto:_FillValue = 1.e+37f;
            rto:long_name="LAPS Fcst storm total precip accum";
            rto:units="m";
            rto:valid_range= 0.f, 1.f;
            rto:LAPS_var="RTO";
            rto:lvl_coord="AGL";
            rto:LAPS_units="M";

        //      LAPS Fcst increment snow accumulation depth
        //      bigfile name = s1hr
        float
            s01(record,z,y,x);
            s01:_FillValue = 1.e+37f;
            s01:long_name="LAPS Fcst increment snow accum depth";
            s01:units="m";
            s01:valid_range= 0.f, 10.f;
            s01:LAPS_var="S01";
            s01:lvl_coord="AGL";
            s01:LAPS_units="M";

        //      LAPS Fcst storm total snow accumulation depth
        //      bigfile name = stot
        float
            sto(record,z,y,x);
            sto:_FillValue = 1.e+37f;
            sto:long_name="LAPS Fcst storm total snow accumulation";
            sto:units="m";
            sto:valid_range= 0.f, 10.f;
            sto:LAPS_var="STO";
            sto:lvl_coord="AGL";
            sto:LAPS_units="M";
	
        //      LAPS Fcst potential temperature   //
        //      not transferred to bigfile
        float
            th(record,z,y,x);
            th:_FillValue = 1.e+37f;
            th:long_name="LAPS Fcst sfc potential temperature";
            th:units="Kelvins";
            th:valid_range= 0.f, 500.f;
            th:LAPS_var="TH";
            th:lvl_coord="AGL";
            th:LAPS_units="K";

        //      LAPS Fcst equivalent potential temperature  //
        //      not transferred to bigfile
        float
            the(record,z,y,x);
            the:_FillValue = 1.e+37f;
            the:long_name="LAPS Fcst sfc equivalent potential temperature";
            the:units="Kelvins";
            the:valid_range= 0.f, 500.f;
            the:LAPS_var="THE";
            the:lvl_coord="AGL";
            the:LAPS_units="K";

        //      LAPS Fcst positive buoyant energy         //
        //      bigfile name = pbe
        float
            pbe(record,z,y,x);
            pbe:_FillValue = 1.e+37f;
            pbe:long_name="LAPS Fcst positive buoyant energy";
            pbe:units="j/kg";
            pbe:valid_range= 0.f, 10000.f;
            pbe:LAPS_var="PBE";
            pbe:lvl_coord="AGL";
            pbe:LAPS_units="J/KG";

         //      LAPS Fcst negative buoyant energy         //
         //      bigfile name = nbe
         float
            nbe(record,z,y,x);
            nbe:_FillValue = 1.e+37f;
            nbe:long_name="LAPS Fcst negative buoyant energy";
            nbe:units="j/kg";
            nbe:valid_range= 0.f, 1000.f;
            nbe:LAPS_var="NBE";
            nbe:lvl_coord="AGL";
            nbe:LAPS_units="J/KG";

        //      LAPS Fcst cloud cover
        //      bigfile name = ccov
        //      not computed yet
        float
            lcv(record,z,y,x);
            lcv:_FillValue = 1.e+37f;
            lcv:long_name="LAPS Fcst cloud cover";
            lcv:units="none";
            lcv:valid_range= 0.f, 1.f;
            lcv:LAPS_var="LCV";
            lcv:lvl_coord="MSL";
            lcv:LAPS_units="FRACTION";

        //      LAPS Fcst cloud ceiling           //
        //      not yet computed -- this is a placeholder
        float
            cce(record,z,y,x);
            cce:_FillValue = 1.e+37f;
            cce:long_name="LAPS Fcst cloud ceiling";
            cce:units="meters";
            cce:valid_range= 0.f, 100000.f;
            cce:LAPS_var="CCE";
            cce:lvl_coord="AGL";
            cce:LAPS_units="M";

        //       LAPS Fcst radar echo tops
        //       bigfile name = mret
        float
            lmt(record,z,y,x);
            lmt:_FillValue = 1.e+37f;
            lmt:long_name="LAPS Fcst radar echo tops";
            lmt:units="meters";
            lmt:valid_range= 0.f, 100000.f;
            lmt:LAPS_var="LMT";
            lmt:lvl_coord="MSL";
            lmt:LAPS_units="M";

        //       LAPS Fcst column max reflectivity
        //       bigfile name = cxr
        float
            lmr(record,z,y,x);
            lmr:_FillValue = 1.e+37f;
            lmr:long_name="LAPS Fcst column max refl";
            lmr:units="dBZ";
            lmr:valid_range= -20.f, 100.f;
            lmr:LAPS_var="LMR";
            lmr:lvl_coord="MSL";
            lmr:LAPS_units="DBZ";

        //       LAPS Fcst low level reflectivity
        //       bigfile name = llr
        float
            llr(record,z,y,x);
            llr:_FillValue = 1.e+37f;
            llr:long_name="LAPS Fcst low level refl";
            llr:units="dBZ";
            llr:valid_range= -20.f, 100.f;
            llr:LAPS_var="LLR";
            llr:lvl_coord="MSL";
            llr:LAPS_units="DBZ";

        //      LAPS Fcst sfc precip type (coded) //
        //      bigfile name = spt
        float
            spt(record,z,y,x);
            spt:_FillValue = 1.e+37f;
            spt:long_name="LAPS Fcst sfc precip type";
            spt:units="code";
            spt:valid_range= 0.f, 100.f;
            spt:LAPS_var="SPT";
            spt:lvl_coord="AGL";
            spt:LAPS_units="CODE";

        //      LAPS Fcst helicity
        //      not transferred to bigfile
        float
            lhe(record,z,y,x);
            lhe:_FillValue = 1.e+37f;
            lhe:long_name="LAPS Fcst helicity";
            lhe:units="m/s**2";
            lhe:valid_range= 0.f, 10000.f;
            lhe:LAPS_var="LHE";
            lhe:lvl_coord="MSL ";
            lhe:LAPS_units="M/S**2";

        //     LAPS Fcst lifted index            //
        //     bigfile name = sli
        float
            li(record,z,y,x);
            li:_FillValue = 1.e+37f;
            li:long_name="LAPS Fcst lifted index";
            li:units="Kelvins";
            li:valid_range= -50.f, 50.f;
            li:LAPS_var="LI";
            li:lvl_coord="AGL";
            li:LAPS_units="K";

         //      LAPS Fcst heat index                      //
         //      bigfile name = hidx
         float
            hi(record,z,y,x);
            hi:_FillValue = 1.e+37f;
            hi:long_name="LAPS Fcst heat index";
            hi:units="Kelvins";
            hi:valid_range= 0.f, 500.f;
            hi:LAPS_var="HI";
            hi:lvl_coord="AGL";
            hi:LAPS_units="K";

         //      LAPS Fcst visibility              //
         //      not computed yet -- this is a placeholder
         float
            vis(record,z,y,x);
            vis:_FillValue = 1.e+37f;
            vis:long_name="LAPS Fcst visibility";
            vis:units="meters";
            vis:valid_range= 0.f, 100000.f;
            vis:LAPS_var="VIS";
            vis:lvl_coord="AGL";
            vis:LAPS_units="M";

        //  	LAPS fire index                     //
        //      bigfile name = fd
        float
            fd(record,z,y,x);
            fd:_FillValue = 1.e+37f;
            fd:long_name="fire index";
            fd:units="none";
            fd:valid_range= 0.f, 20.f;
            fd:LAPS_var="FD";
            fd:lvl_coord="AGL";
            fd:LAPS_units="NONE";

        //      Model Topography                    //
        //      bigfile name = 
        float
            ter(record,z,y,x);
            ter:_FillValue = 1.e+37f;
            ter:long_name="terrain height";
            ter:units="meters";
            ter:valid_range= -200.f, 20000.f;
            ter:LAPS_var="TER";
            ter:lvl_coord="MSL";
            ter:LAPS_units="METERS";           

        //	LAPS variables
                	        
        long
            imax,
            jmax,
            kmax,
            kdim;

        char
            u_comment(record,z,namelen),
            v_comment(record,z,namelen),
            w_comment(record,z,namelen),
            t_comment(record,z,namelen),
            td_comment(record,z,namelen),
            rh_comment(record,z,namelen),
            lcb_comment(record,z,namelen),
            lct_comment(record,z,namelen),
            msl_comment(record,z,namelen),
            p_comment(record,z,namelen),
            ps_comment(record,z,namelen),
            lil_comment(record,z,namelen),
            tpw_comment(record,z,namelen),
            r01_comment(record,z,namelen),
            rto_comment(record,z,namelen),
            s01_comment(record,z,namelen),
            sto_comment(record,z,namelen),
            th_comment(record,z,namelen),
            the_comment(record,z,namelen),
            pbe_comment(record,z,namelen),
            nbe_comment(record,z,namelen),
            lcv_comment(record,z,namelen),
            cce_comment(record,z,namelen),
            lmt_comment(record,z,namelen),
            lmr_comment(record,z,namelen),
            llr_comment(record,z,namelen),
            spt_comment(record,z,namelen),
            lhe_comment(record,z,namelen),
            li_comment(record,z,namelen),
            hi_comment(record,z,namelen),
            vis_comment(record,z,namelen),
            fd_comment(record,z,namelen),
            ter_comment(record,z.namelen),
            asctime(record,namelen);

			
        //	inventory variables

        short
            u_fcinv(record, z);
            u_fcinv:_FillValue= 0s;
              	
        short
            v_fcinv(record, z);
            v_fcinv:_FillValue= 0s;
              	
        short
            w_fcinv(record, z);
            w_fcinv:_FillValue= 0s;
              	
        short
            t_fcinv(record, z);
            t_fcinv:_FillValue= 0s;
              	
        short
            td_fcinv(record, z);
            td_fcinv:_FillValue= 0s;
              	
        short
            rh_fcinv(record, z);
            rh_fcinv:_FillValue= 0s;

        short
            lcb_fcinv(record, z);
            lcb_fcinv:_FillValue= 0s;

        short
            lct_fcinv(record, z);
            lct_fcinv:_FillValue= 0s;

        short
            msl_fcinv(record, z);
            msl_fcinv:_FillValue= 0s;

        short
            p_fcinv(record, z);
            p_fcinv:_FillValue= 0s;
              	
        short
            ps_fcinv(record, z);
            ps_fcinv:_FillValue= 0s;

        short
            lil_fcinv(record, z);
            lil_fcinv:_FillValue= 0s;

        short
            tpw_fcinv(record, z);
            tpw_fcinv:_FillValue= 0s;

        short
            r01_fcinv(record, z);
            r01_fcinv:_FillValue= 0s;

        short
            rto_fcinv(record, z);
            rto_fcinv:_FillValue= 0s;

        short
            s01_fcinv(record, z);
            s01_fcinv:_FillValue= 0s;

        short
            sto_fcinv(record, z);
            sto_fcinv:_FillValue= 0s;

        short
            th_fcinv(record, z);
            th_fcinv:_FillValue= 0s;

        short
            the_fcinv(record, z);
            the_fcinv:_FillValue= 0s;

        short
            pbe_fcinv(record, z);
            pbe_fcinv:_FillValue= 0s;

        short
            nbe_fcinv(record, z);
            nbe_fcinv:_FillValue= 0s;

        short
            lcv_fcinv(record, z);
            lcv_fcinv:_FillValue= 0s;

        short
            cce_fcinv(record, z);
            cce_fcinv:_FillValue= 0s;

        short
            lmt_fcinv(record, z);
            lmt_fcinv:_FillValue= 0s;

        short
            lmr_fcinv(record, z);
            lmr_fcinv:_FillValue= 0s;

        short
            llr_fcinv(record, z);
            llr_fcinv:_FillValue= 0s;

        short
            spt_fcinv(record, z);
            spt_fcinv:_FillValue= 0s;

        short
            lhe_fcinv(record, z);
            lhe_fcinv:_FillValue= 0s;

        short
            li_fcinv(record, z);
            li_fcinv:_FillValue= 0s;

        short
            hi_fcinv(record, z);
            hi_fcinv:_FillValue= 0s;

        short
            vis_fcinv(record, z);
            vis_fcinv:_FillValue= 0s;

        short
            fd_fcinv(record, z);
            fd_fcinv:_FillValue= 0s;

        short
            ter_fcinv(record, z);
            ter_fcinv:_FillValue= 0s;   

        //	list of grid levels

        float 
            level(z);
            level:long_name="level of data";
	    level:units = "hectopascals";
                    	
        //      validtime of the grid 

        double
            valtime(record);
            valtime:long_name = "valid time";
            valtime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      reference time of the process

        double
            reftime(record);
            reftime:long_name = "reference time";
            reftime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      nice name for originating center

        char
            origin_name(namelen);

        //      nice name for process

        char
            process_name(namelen);

        //      nice name for grid description instance
        char
            grid_name(namelen);

        //      basic assumption about earth shape
        char
            earth_shape(namelen);

        // navigation variables using 
        // WMO FM 92-VIII Ext.GRIB specification names
  
        char    grid_type(nav, namelen);
                grid_type:long_name = "GRIB-1 grid type";
  
        char    x_dim(nav, namelen);
                x_dim:long_name = "longitude dimension";
  
        char    y_dim(nav, namelen);
                y_dim:long_name = "latitude dimension";
  
        short   Nx(nav);
                Nx:long_name = "number of x points";
  
        short   Ny(nav);
                Ny:long_name =  "number of y points";
  
        float   La1(nav);
                La1:long_name = "first latitude";
                La1:units = "degrees_north";
  
        float   Lo1(nav);
                Lo1:long_name = "first longitude";
                Lo1:units = "degrees_east" ;
    
        float   LoV(nav);
                LoV:long_name = "orientation of grid" ;
                LoV:units = "degrees_east";
  
        float   Latin1(nav);
                Latin1:long_name = "orientation of grid" ;
                Latin1:units = "degrees_north";

        float   Latin2(nav);
                Latin2:long_name = "orientation of grid" ;
                Latin2:units = "degrees_north";

        float   Dx(nav);
                Dx:long_name = "x grid increment";
                Dx:units = "kilometers";
  
        float   Dy(nav);
                Dy:long_name = "y grid increment";
                Dy:units = "kilometers";
  
        // end of navigation variables

        :Conventions = "NUWG";
        :history = "created by LAPS Branch of FSL";
        :record = "valtime, reftime";
        :title = "LAPS rsf file - forecast model surface data";
        :version = 3;

    data:

        earth_shape     = "spherical radius";
        grid_name       = "LAPS rsf file - forecast model surface data";
        process_name    = "LAPS - Local Analysis and Prediction System";
        x_dim           = "x";
        y_dim           = "y";
}                       
