netcdf lsx {

    dimensions:
        record = unlimited,
        z = 1,
	x = 125,
	y = 105,
        nav = 1,
        namelen = 132;
		
    variables:
        //	surface u wind component

	float                                  
            u(record,z,y,x);
            u:navigation_dim = "nav";
            u:record = "valtime, reftime";
            u:_FillValue = 1.e+37f;
            u:long_name="u-component of surface wind";
            u:units="meters / second";
            u:valid_range= -200.f, 200.f;
            u:LAPS_var="U";
            u:lvl_coord="AGL";
	    u:LAPS_units="M/S";

        //      surface v wind component        //

        float
            v(record,z,y,x);
            v:long_name="v-component of surface wind";
            v:navigation_dim = "nav";
            v:record = "valtime, reftime";
            v:_FillValue = 1.e+37f;
            v:units="meters/second";
            v:valid_range= -200.f, 200.f;
            v:LAPS_var="V";
            v:lvl_coord="AGL";
            v:LAPS_units="M/S";
 
        //      1500 M Reduced Pressure         //

        float
            p(record,z,y,x);
            p:navigation_dim = "nav";
            p:record = "valtime, reftime";
            p:_FillValue = 1.e+37f;
            p:long_name="1500 m reduced pressure";
            p:units="pascals";
            p:valid_range= 0.f, 1000.f;
            p:LAPS_var="P";
            p:lvl_coord="AGL ";
            p:LAPS_units="PA";
 
        //      surface temperature     //

        float
            t(record,z,y,x);
            t:navigation_dim = "nav";
            t:record = "valtime, reftime";
            t:_FillValue = 1.e+37f;
            t:long_name="surface temperature";
            t:units="degrees kelvin";
            t:valid_range= -150.f, 150.f;
            t:LAPS_var="T";
            t:lvl_coord="AGL ";
            t:LAPS_units="K";

        //      surface dewpoint temperature    //

        float
            td(record,z,y,x);
            td:navigation_dim = "nav";
            td:record = "valtime, reftime";
            td:_FillValue = 1.e+37f;
            td:long_name="surface dewpoint temperature";
            td:units="degrees kelvin";
            td:valid_range= -75.f, 125.f;
            td:LAPS_var="TD";
            td:lvl_coord="AGL ";
            td:LAPS_units="K";
 
        //      Vertical Velocity       //

        float
            vv(record,z,y,x);
            vv:navigation_dim = "nav";
            vv:record = "valtime, reftime";
            vv:_FillValue = 1.e+37f;
            vv:long_name="vertical velocity";
            vv:units="meters/second";
            vv:valid_range= 0.f, 20000.f;
            vv:LAPS_var="VV";
            vv:lvl_coord="AGL";
            vv:LAPS_units="M/S";

        //      Relative humidity       //

        float
            rh(record,z,y,x);
            rh:navigation_dim = "nav";
            rh:record = "valtime, reftime";
            rh:_FillValue = 1.e+37f;
            rh:long_name="relative humidity";
            rh:units="meters";
            rh:valid_range= -20000.f, 20000.f;
            rh:LAPS_var="RH";
            rh:lvl_coord="AGL";
            rh:LAPS_units="M";

        //      MSL Pressure            //

        float
            msl(record,z,y,x);
            msl:navigation_dim = "nav";
            msl:record = "valtime, reftime";
            msl:_FillValue = 1.e+37f;
            msl:long_name="MSL pressure";
            msl:units="pascals";
            msl:valid_range= -20000.f, 20000.f;
            msl:LAPS_var="MSL";
            msl:lvl_coord="AGL";
            msl:LAPS_units="PA";
 
        //      Temperature Advection   //

        float
            tad(record,z,y,x);
            tad:navigation_dim = "nav";
            tad:record = "valtime, reftime";
            tad:_FillValue = 1.e+37f;
            tad:long_name="temperature advection";
            tad:units="degrees Kelvin/second";
            tad:valid_range= -20000.f, 20000.f;
            tad:LAPS_var="TAD";
            tad:lvl_coord="MSL";
            tad:LAPS_units="K/S";
 
        //      Potential temperature   //

        float
            th(record,z,y,x);
            th:navigation_dim = "nav";
            th:record = "valtime, reftime";
            th:_FillValue = 1.e+37f;
            th:long_name="potential temperature";
            th:units="degrees Kelvin";
            th:valid_range= -75.f, 125.f;
            th:LAPS_var="TH";
            th:lvl_coord="AGL";
            th:LAPS_units="K";
 
        //      equivalent potential temperature  //

        float
            the(record,z,y,x);
            the:navigation_dim = "nav";
            the:record = "valtime, reftime";
            the:_FillValue = 1.e+37f;
            the:long_name="equivalent potential temperature";
            the:units="degrees Kelvin";
            the:valid_range= -20000.f, 20000.f;
            the:LAPS_var="THE";
            the:lvl_coord="AGL";
            the:LAPS_units="K";
 
        //      surface pressure        //

        float
            ps(record,z,y,x);
            ps:navigation_dim = "nav";
            ps:record = "valtime, reftime";
            ps:_FillValue = 1.e+37f;
            ps:long_name="surface pressure";
            ps:units="pascals";
            ps:valid_range= -20000.f, 20000.f;
            ps:LAPS_var="PS";
            ps:lvl_coord="AGL";
            ps:LAPS_units="PA";
 
        //      vorticity               //

        float
            vor(record,z,y,x);
            vor:navigation_dim = "nav";
            vor:record = "valtime, reftime";
            vor:_FillValue = 1.e+37f;
            vor:long_name="vorticity";
            vor:units="/second";
            vor:valid_range= -20000.f, 20000.f;
            vor:LAPS_var="VOR";
            vor:lvl_coord="AGL";
            vor:LAPS_units="/S";

        //      mixing ratio            //

        float
            mr(record,z,y,x);
            mr:navigation_dim = "nav";
            mr:record = "valtime, reftime";
            mr:_FillValue = 1.e+37f;
            mr:long_name="mixing ratio";
            mr:units="grams/kikogram";
            mr:valid_range= -20000.f, 20000.f;
            mr:LAPS_var="MR";
            mr:lvl_coord="AGL";
            mr:LAPS_units="G/KG";
 
        //      moisture convergence            //

        float
            mrc(record,z,y,x);
            mrc:navigation_dim = "nav";
            mrc:record = "valtime, reftime";
            mrc:_FillValue = 1.e+37f;
            mrc:long_name="moisture convergence";
            mrc:units="grams/kilogram/seconds";
            mrc:valid_range= -20000.f, 20000.f;
            mrc:LAPS_var="MRC";
            mrc:lvl_coord="AGL";
            mrc:LAPS_units="G/KG/S";
 
        //      divergence              //

        float
            div(record,z,y,x);
            div:navigation_dim = "nav";
            div:record = "valtime, reftime";
            div:_FillValue = 1.e+37f;
            div:long_name="divergence";
            div:units="/second";
            div:valid_range= -20000.f, 20000.f;
            div:LAPS_var="DIV";
            div:lvl_coord="AGL";
            div:LAPS_units="/S";
 
        //      potential temperature advection         //

        float
            tha(record,z,y,x);
            tha:navigation_dim = "nav";
            tha:record = "valtime, reftime";
            tha:_FillValue = 1.e+37f;
            tha:long_name="potential temperature advection";
            tha:units="kilograms/second";
            tha:valid_range= -20000.f, 20000.f;
            tha:LAPS_var="THA";
            tha:lvl_coord="AGL";
            tha:LAPS_units="K/S";
 
        //      moisture advection      //

        float
            mra(record,z,y,x);
            mra:navigation_dim = "nav";
            mra:record = "valtime, reftime";
            mra:_FillValue = 1.e+37f;
            mra:long_name="moisture advection";
            mra:units="grams/kilogram/second";
            mra:valid_range= -20000.f, 20000.f;
            mra:LAPS_var="MRA";
            mra:lvl_coord="AGL";
            mra:LAPS_units="G/KG/S";
 
        //      surface wind speed      //
        float
            spd(record,z,y,x);
            spd:navigation_dim = "nav";
            spd:record = "valtime, reftime";
            spd:_FillValue = 1.e+37f;
            spd:long_name="surface wind speed";
            spd:units="meters/second";
            spd:valid_range= -20000.f, 20000.f;
            spd:LAPS_var="SPD";
            spd:lvl_coord="AGL";
            spd:LAPS_units="M/S";
 
        //      colorado severe storm index     //

        float
            css(record,z,y,x);
            css:navigation_dim = "nav";
            css:record = "valtime, reftime";
            css:_FillValue = 1.e+37f;
            css:long_name="colorado severe storm index";
            css:units="          ";
            css:valid_range= -20000.f, 20000.f;
            css:LAPS_var="CSS";
            css:lvl_coord="AGL";
            css:LAPS_units="          ";
 
         //      visability              //

         float
            vis(record,z,y,x);
            vis:navigation_dim = "nav";
            vis:record = "valtime, reftime";
            vis:_FillValue = 1.e+37f;
            vis:long_name="visibility";
            vis:units="meters";
            vis:valid_range= -20000.f, 20000.f;
            vis:LAPS_var="VIS";
            vis:lvl_coord="AGL";
            vis:LAPS_units="M";
 
         //      fire weather index              //
         float
            fwx(record,z,y,x);
            fwx:navigation_dim = "nav";
            fwx:record = "valtime, reftime";
            fwx:_FillValue = 1.e+37f;
            fwx:long_name="Fire danger";
            fwx:units="none";
            fwx:valid_range= 0.f, 20.f;
            fwx:LAPS_var="FWX";
            fwx:lvl_coord="none";
            fwx:LAPS_units="none";
 
         //      heat index                      //
         float
            hi(record,z,y,x);
            hi:navigation_dim = "nav";
            hi:record = "valtime, reftime";
            hi:_FillValue = 1.e+37f;
            hi:long_name="Heat index";
            hi:units="none";
            hi:valid_range= 0.f, 20.f;
            hi:LAPS_var="HI";
            hi:lvl_coord="none";
            hi:LAPS_units="none";

        //      ground temperature
        float
            tgd(record,z,y,x);
            tgd:_FillValue = 1.e+37f;
            tgd:long_name="Ground Temperature";
            tgd:units="K";
            tgd:valid_range= 0.f, 400.f;
            tgd:LAPS_var="TGD";
            tgd:lvl_coord="AGL";
            tgd:LAPS_units="K";

                	        
        //	LAPS variables

        long
            imax,
            jmax,
            kmax,
            kdim;

        char
            u_comment(record,z,namelen),
            v_comment(record,z,namelen),
            p_comment(record,z,namelen),
            t_comment(record,z,namelen),
            td_comment(record,z,namelen),
            vv_comment(record,z,namelen),
            rh_comment(record,z,namelen),
            msl_comment(record,z,namelen),
            tad_comment(record,z,namelen),
            th_comment(record,z,namelen),
            the_comment(record,z,namelen),
            ps_comment(record,z,namelen),
            vor_comment(record,z,namelen),
            mr_comment(record,z,namelen),
            mrc_comment(record,z,namelen),
            div_comment(record,z,namelen),
            tha_comment(record,z,namelen),
            mra_comment(record,z,namelen),
            spd_comment(record,z,namelen),
            css_comment(record,z,namelen),
            vis_comment(record,z,namelen),
            fwx_comment(record,z,namelen),
            hi_comment(record,z,namelen),
            tgd_comment(record,z,namelen),
            asctime(record,namelen);

			
        //	inventory variables

        short
            u_fcinv(record, z);
            u_fcinv:_FillValue= 0s;
              	
        short
            v_fcinv(record, z);
            v_fcinv:_FillValue= 0s;
              	
        short
            p_fcinv(record, z);
            p_fcinv:_FillValue= 0s;
              	
        short
            t_fcinv(record, z);
            t_fcinv:_FillValue= 0s;
              	
        short
            td_fcinv(record, z);
            td_fcinv:_FillValue= 0s;
              	
        short
            vv_fcinv(record, z);
            vv_fcinv:_FillValue= 0s;
              	
        short
            rh_fcinv(record, z);
            rh_fcinv:_FillValue= 0s;
              	
        short
            msl_fcinv(record, z);
            msl_fcinv:_FillValue= 0s;
              	
        short
            tad_fcinv(record, z);
            tad_fcinv:_FillValue= 0s;
              	
        short
            th_fcinv(record, z);
            th_fcinv:_FillValue= 0s;
              	
        short
            the_fcinv(record, z);
            the_fcinv:_FillValue= 0s;
              	
        short
            ps_fcinv(record, z);
            ps_fcinv:_FillValue= 0s;
              	
        short
            vor_fcinv(record, z);
            vor_fcinv:_FillValue= 0s;
              	
        short
            mr_fcinv(record, z);
            mr_fcinv:_FillValue= 0s;
              	
        short
            mrc_fcinv(record, z);
            mrc_fcinv:_FillValue= 0s;
              	
        short
            div_fcinv(record, z);
            div_fcinv:_FillValue= 0s;
              	
        short
            tha_fcinv(record, z);
            tha_fcinv:_FillValue= 0s;
              	
        short
            mra_fcinv(record, z);
            mra_fcinv:_FillValue= 0s;
              	
        short
            spd_fcinv(record, z);
            spd_fcinv:_FillValue= 0s;
              	
        short
            css_fcinv(record, z);
            css_fcinv:_FillValue= 0s;
              	
        short
            vis_fcinv(record, z);
            vis_fcinv:_FillValue= 0s;
              	
        short
            fwx_fcinv(record, z);
            fwx_fcinv:_FillValue= 0s;
              	
        short
            hi_fcinv(record, z);
            hi_fcinv:_FillValue= 0s;
              	
        short
            tgd_fcinv(record, z);
            tgd_fcinv:_FillValue= 0s;
              	
        //	list of grid levels

        float 
            level(z);
            level:long_name="level of data";
	    level:units = "hectopascals";
                    	
        //      validtime of the grid 

        double
            valtime(record);
            valtime:long_name = "valid time";
            valtime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      reference time of the process

        double
            reftime(record);
            reftime:long_name = "reference time";
            reftime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      nice name for originating center

        char
            origin_name(namelen);

        //      nice name for process

        char
            process_name(namelen);

        //      nice name for grid description instance
        char
            grid_name(namelen);

        //      basic assumption about earth shape
        char
            earth_shape(namelen);

        // navigation variables using 
        // WMO FM 92-VIII Ext.GRIB specification names
  
        char    grid_type(nav, namelen);
                grid_type:long_name = "GRIB-1 grid type";
  
        char    x_dim(nav, namelen);
                x_dim:long_name = "longitude dimension";
  
        char    y_dim(nav, namelen);
                y_dim:long_name = "latitude dimension";
  
        short   Nx(nav);
                Nx:long_name = "number of x points";
  
        short   Ny(nav);
                Ny:long_name =  "number of y points";
  
        float   La1(nav);
                La1:long_name = "first latitude";
                La1:units = "degrees_north";
  
        float   Lo1(nav);
                Lo1:long_name = "first longitude";
                Lo1:units = "degrees_east" ;
    
        float   LoV(nav);
                LoV:long_name = "orientation of grid" ;
                LoV:units = "degrees_east";
  
        float   Latin1(nav);
                Latin1:long_name = "orientation of grid" ;
                Latin1:units = "degrees_north";

        float   Latin2(nav);
                Latin2:long_name = "orientation of grid" ;
                Latin2:units = "degrees_north";

        float   Dx(nav);
                Dx:long_name = "x grid increment";
                Dx:units = "kilometers";
  
        float   Dy(nav);
                Dy:long_name = "y grid increment";
                Dy:units = "kilometers";
  
        // end of navigation variables

        :Conventions = "NUWG";
        :history = "created by LAPS Branch of FSL";
        :record = "valtime, reftime";
        :title = "LAPS lsx file - LAPS surface";
        :version = 3;

    data:

        earth_shape     = "spherical radius";
        grid_name       = "LAPS lsx file - LAPS surface";
        process_name    = "LAPS - Local Analysis and Prediction System";
        x_dim           = "x";
        y_dim           = "y";
}                       
