netcdf rsf {

    dimensions:
        record = unlimited,
        z = 1,
	x = 61,
	y = 61,
        nav = 1,
        namelen = 132;
		
    variables:

        //	LAPS Fcst sfc u wind component
	float                                  
            u(record,z,y,x);
            u:_FillValue = 1.e+37f;
            u:long_name="LAPS Fcst sfc u wind component";
            u:units="m/s";
            u:valid_range= -200.f, 200.f;
            u:LAPS_var="U";
            u:lvl_coord="AGL";
	    u:LAPS_units="M/S";
                	        
        //	LAPS Fcst sfc v wind component
	float                                  
            v(record,z,y,x);
            v:_FillValue = 1.e+37f;
            v:long_name="LAPS Fcst sfc v wind component";
            v:units="m/s";
            v:valid_range= -200.f, 200.f;
            v:LAPS_var="V";
            v:lvl_coord="AGL";
	    v:LAPS_units="M/S";
                	        
                	        
        //	LAPS Fcst sfc temperature
	float                                  
            t(record,z,y,x);
            t:_FillValue = 1.e+37f;
            t:long_name="LAPS Fcst sfc temperature";
            t:units="Kelvins";
            t:valid_range= 0.f, 500.f;
            t:LAPS_var="T";
            t:lvl_coord="AGL";
	    t:LAPS_units="K";
                	        
        //	LAPS Fcst surface dewpoint
	float                                  
            td(record,z,y,x);
            td:_FillValue = 1.e+37f;
            td:long_name="LAPS Fcst sfc dewpoint";
            td:units="Kelvins";
            td:valid_range= 0.f, 500.f;
            td:LAPS_var="TD";
            td:lvl_coord="AGL";
	    td:LAPS_units="K";

        //      LAPS Fcst relative humidity       //
        //      bigfile name = rh
        float
            rh(record,z,y,x);
            rh:_FillValue = 1.e+37f;
            rh:long_name="LAPS Fcst sfc relative humidity";
            rh:units="meters";
            rh:valid_range= 0.f, 100.f;
            rh:LAPS_var="RH";
            rh:lvl_coord="AGL";
            rh:LAPS_units="PERCENT";

        //      LAPS Fcst MSL Pressure            //
        //      bigfile name = mslp
        float
            msl(record,z,y,x);
            msl:_FillValue = 1.e+37f;
            msl:long_name="LAPS Fcst MSL pressure";
            msl:units="pascals";
            msl:valid_range= 0.f, 100000.f;
            msl:LAPS_var="MSL";
            msl:lvl_coord="MSL";
            msl:LAPS_units="PA";

                	        
        //      LAPS Fcst surface pressure (looks like topo)      //

        float
            ps(record,z,y,x);
            ps:_FillValue = 1.e+37f;
            ps:long_name="LAPS Fcst sfc pressure";
            ps:units="pascals";
            ps:valid_range= 0.f, 100000.f;
            ps:LAPS_var="PS";
            ps:lvl_coord="AGL";
            ps:LAPS_units="PA";

        //      LAPS Fcst potential temperature   //
        float
            th(record,z,y,x);
            th:_FillValue = 1.e+37f;
            th:long_name="LAPS Fcst sfc potential temperature";
            th:units="Kelvins";
            th:valid_range= 0.f, 500.f;
            th:LAPS_var="TH";
            th:lvl_coord="AGL";
            th:LAPS_units="K";

        //      LAPS Fcst equivalent potential temperature  //
        float
            the(record,z,y,x);
            the:_FillValue = 1.e+37f;
            the:long_name="LAPS Fcst sfc equivalent potential temperature";
            the:units="Kelvins";
            the:valid_range= 0.f, 500.f;
            the:LAPS_var="THE";
            the:lvl_coord="AGL";
            the:LAPS_units="K";



        //	LAPS variables
                	        
        long
            imax,
            jmax,
            kmax,
            kdim;

        char
            u_comment(record,z,namelen),
            v_comment(record,z,namelen),
            t_comment(record,z,namelen),
            rh_comment(record,z,namelen),
            td_comment(record,z,namelen),
            msl_comment(record,z,namelen),
            ps_comment(record,z,namelen),
            th_comment(record,z,namelen),
            the_comment(record,z,namelen),
            asctime(record,namelen);

			
        //	inventory variables

        short
            u_fcinv(record, z);
            u_fcinv:_FillValue= 0s;
              	
        short
            v_fcinv(record, z);
            v_fcinv:_FillValue= 0s;
              	
        short
            t_fcinv(record, z);
            t_fcinv:_FillValue= 0s;
              	
        short
            td_fcinv(record, z);
            td_fcinv:_FillValue= 0s;
              	
        short
            rh_fcinv(record, z);
            rh_fcinv:_FillValue= 0s;

        short
            msl_fcinv(record, z);
            msl_fcinv:_FillValue= 0s;

        short
            ps_fcinv(record, z);
            ps_fcinv:_FillValue= 0s;

        short
            th_fcinv(record, z);
            th_fcinv:_FillValue= 0s;

        short
            the_fcinv(record, z);
            the_fcinv:_FillValue= 0s;

        //	list of grid levels

        float 
            level(z);
            level:long_name="level of data";
	    level:units = "hectopascals";
                    	
        //      validtime of the grid 

        double
            valtime(record);
            valtime:long_name = "valid time";
            valtime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      reference time of the process

        double
            reftime(record);
            reftime:long_name = "reference time";
            reftime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      nice name for originating center

        char
            origin_name(namelen);

        //      nice name for process

        char
            process_name(namelen);

        //      nice name for grid description instance
        char
            grid_name(namelen);

        //      basic assumption about earth shape
        char
            earth_shape(namelen);

        // navigation variables using 
        // WMO FM 92-VIII Ext.GRIB specification names
  
        char    grid_type(nav, namelen);
                grid_type:long_name = "GRIB-1 grid type";
  
        char    x_dim(nav, namelen);
                x_dim:long_name = "longitude dimension";
  
        char    y_dim(nav, namelen);
                y_dim:long_name = "latitude dimension";
  
        short   Nx(nav);
                Nx:long_name = "number of x points";
  
        short   Ny(nav);
                Ny:long_name =  "number of y points";
  
        float   La1(nav);
                La1:long_name = "first latitude";
                La1:units = "degrees_north";
  
        float   Lo1(nav);
                Lo1:long_name = "first longitude";
                Lo1:units = "degrees_east" ;
    
        float   LoV(nav);
                LoV:long_name = "orientation of grid" ;
                LoV:units = "degrees_east";
  
        float   Latin1(nav);
                Latin1:long_name = "orientation of grid" ;
                Latin1:units = "degrees_north";

        float   Latin2(nav);
                Latin2:long_name = "orientation of grid" ;
                Latin2:units = "degrees_north";

        float   Dx(nav);
                Dx:long_name = "x grid increment";
                Dx:units = "kilometers";
  
        float   Dy(nav);
                Dy:long_name = "y grid increment";
                Dy:units = "kilometers";
  
        // end of navigation variables

        :Conventions = "NUWG";
        :history = "created by LAPS Branch of FSL";
        :record = "valtime, reftime";
        :title = "LAPS rsf file - forecast model surface data";
        :version = 3;

    data:

        earth_shape     = "spherical radius";
        grid_name       = "LAPS rsf file - forecast model surface data";
        process_name    = "LAPS - Local Analysis and Prediction System";
        x_dim           = "x";
        y_dim           = "y";
}                       
