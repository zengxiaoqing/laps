netcdf rsf {

    dimensions:
        record = unlimited,
        z = 1,
	x = 125,
	y = 105,
        nav = 1,
        namelen = 132;
		
    variables:
        //	LAPS Fcst sfc wind component

	float                                  
            u(record,z,y,x);
            u:navigation_dim = "nav";
            u:record = "valtime, reftime";
            u:_FillValue = 1.e+37f;
            u:long_name="LAPS Fcst sfc u wind component";
            u:units="meters / second";
            u:valid_range= -200.f, 200.f;
            u:LAPS_var="U";
            u:lvl_coord="HPA";
	    u:LAPS_units="M/S";
                	        
        //	LAPS Fcst sfc v wind component

	float                                  
            v(record,z,y,x);
            v:navigation_dim = "nav";
            v:record = "valtime, reftime";
            v:_FillValue = 1.e+37f;
            v:long_name="LAPS Fcst sfc v wind component";
            v:units="meters / second";
            v:valid_range= -200.f, 200.f;
            v:LAPS_var="V";
            v:lvl_coord="HPA";
	    v:LAPS_units="M/S";
                	        
        //	LAPS Fcst sfc temperature

	float                                  
            t(record,z,y,x);
            t:navigation_dim = "nav";
            t:record = "valtime, reftime";
            t:_FillValue = 1.e+37f;
            t:long_name="LAPS Fcst surface temperature";
            t:units="degrees Kelvin";
            t:valid_range= -200.f, 200.f;
            t:LAPS_var="T";
            t:lvl_coord="AGL";
	    t:LAPS_units="K";
                	        
        //	LAPS Fcst 1500m pressure

	float                                  
            p(record,z,y,x);
            p:navigation_dim = "nav";
            p:record = "valtime, reftime";
            p:_FillValue = 1.e+37f;
            p:long_name="LAPS Fcst 1500m pressure";
            p:units="pascals";
            p:valid_range= -200.f, 200.f;
            p:LAPS_var="P";
            p:lvl_coord="AGL";
	    p:LAPS_units="PA";
                	        
        //	LAPS Fcst surface dewpoint

	float                                  
            td(record,z,y,x);
            td:navigation_dim = "nav";
            td:record = "valtime, reftime";
            td:_FillValue = 1.e+37f;
            td:long_name="LAPS Fcst surface dewpoint";
            td:units="degrees Kelvin";
            td:valid_range= -200.f, 200.f;
            td:LAPS_var="TD";
            td:lvl_coord="AGL";
	    td:LAPS_units="K";

        //      Relative humidity       //

        float
            rh(record,z,y,x);
            rh:navigation_dim = "nav";
            rh:record = "valtime, reftime";
            rh:_FillValue = 1.e+37f;
            rh:long_name="LAPS Fcst relative humidity";
            rh:units="meters";
            rh:valid_range= -20000.f, 20000.f;
            rh:LAPS_var="RH";
            rh:lvl_coord="AGL";
            rh:LAPS_units="M";

        //      cloud base

        float
            lcb(record,z,y,x);
            lcb:navigation_dim = "nav";
            lcb:record = "valtime, reftime";
            lcb:_FillValue = 1.e+37f;
            lcb:long_name="LAPS cloud base";
            lcb:units="meters";
            lcb:valid_range= -200.f, 200.f;
            lcb:LAPS_var="LCB";
            lcb:lvl_coord="MSL";
            lcb:LAPS_units="M";
        //      cloud top

        float
            lct(record,z,y,x);
            lct:navigation_dim = "nav";
            lct:record = "valtime, reftime";
            lct:_FillValue = 1.e+37f;
            lct:long_name="LAPS cloud top";
            lct:units="meters";
            lct:valid_range= -200.f, 200.f;
            lct:LAPS_var="LCT";
            lct:lvl_coord="MSL";
            lct:LAPS_units="M";

        //      MSL Pressure            //

        float
            msl(record,z,y,x);
            msl:navigation_dim = "nav";
            msl:record = "valtime, reftime";
            msl:_FillValue = 1.e+37f;
            msl:long_name="MSL pressure";
            msl:units="pascals";
            msl:valid_range= -20000.f, 20000.f;
            msl:LAPS_var="MSL";
            msl:lvl_coord="AGL";
            msl:LAPS_units="PA";

        //      integrated liquid water

        float
            lil(record,z,y,x);
            lil:navigation_dim = "nav";
            lil:record = "valtime, reftime";
            lil:_FillValue = 1.e+37f;
            lil:long_name="integrated liquid water";
            lil:units="grams/meter**2";
            lil:valid_range= 0.f, 100.f;
            lil:LAPS_var="LIL";
            lil:lvl_coord="MSL";
            lil:LAPS_units="G/M**2";

        //      integrated total precip water

        float
            tpw(record,z,y,x);
            tpw:navigation_dim = "nav";
            tpw:record = "valtime, reftime";
            tpw:_FillValue = 1.e+37f;
            tpw:long_name="integrated total precipitable water";
            tpw:units="meters";
            tpw:valid_range= 0.f, 0.100f;
            tpw:LAPS_var="TPW";
            tpw:lvl_coord="    ";
            tpw:LAPS_units="M";

        //      60 minute precip accumulation

        float
            r01(record,z,y,x);
            r01:navigation_dim = "nav";
            r01:record = "valtime, reftime";
            r01:_FillValue = 1.e+37f;
            r01:long_name="LAPS 60 minute precip. accum.";
            r01:units="meters";
            r01:valid_range= -200.f, 200.f;
            r01:LAPS_var="R01";
            r01:lvl_coord="MSL";
            r01:LAPS_units="M";

        //      storm total precip accum

        float
            rto(record,z,y,x);
            rto:navigation_dim = "nav";
            rto:record = "valtime, reftime";
            rto:_FillValue = 1.e+37f;
            rto:long_name="storm total precip. accum.";
            rto:units="meters";
            rto:valid_range= -200.f, 200.f;
            rto:LAPS_var="RTO";
            rto:lvl_coord="MSL";
            rto:LAPS_units="M";

        //      60 min snow accumulation

        float
            s01(record,z,y,x);
            s01:navigation_dim = "nav";
            s01:record = "valtime, reftime";
            s01:_FillValue = 1.e+37f;
            s01:long_name="LAPS 60 minute snow accum.";
            s01:units="meters";
            s01:valid_range= -200.f, 200.f;
            s01:LAPS_var="S01";
            s01:lvl_coord="MSL";
            s01:LAPS_units="M";

        //      storm total accumulation

        float
            sto(record,z,y,x);
            sto:navigation_dim = "nav";
            sto:record = "valtime, reftime";
            sto:_FillValue = 1.e+37f;
            sto:long_name="storm total snow accumulation";
            sto:units="meters";
            sto:valid_range= -200.f, 200.f;
            sto:LAPS_var="STO";
            sto:lvl_coord="MSL";
            sto:LAPS_units="M";
	
        //      Potential temperature   //

        float
            th(record,z,y,x);
            th:navigation_dim = "nav";
            th:record = "valtime, reftime";
            th:_FillValue = 1.e+37f;
            th:long_name="LAPS Fcst potential temperature";
            th:units="degrees Kelvin";
            th:valid_range= -75.f, 125.f;
            th:LAPS_var="TH";
            th:lvl_coord="AGL";
            th:LAPS_units="K";

        //      equivalent potential temperature  //

        float
            the(record,z,y,x);
            the:navigation_dim = "nav";
            the:record = "valtime, reftime";
            the:_FillValue = 1.e+37f;
            the:long_name="LAPS Fcst equivalent potential temperature";
            the:units="degrees Kelvin";
            the:valid_range= -20000.f, 20000.f;
            the:LAPS_var="THE";
            the:lvl_coord="AGL";
            the:LAPS_units="K";

        //      positive buoyant energy         //
        float
            pbe(record,z,y,x);
            pbe:navigation_dim = "nav";
            pbe:record = "valtime, reftime";
            pbe:_FillValue = 1.e+37f;
            pbe:long_name="positive buoyant energy";
            pbe:units="joules/kilogram";
            pbe:valid_range= -20000.f, 20000.f;
            pbe:LAPS_var="PBE";
            pbe:lvl_coord="AGL";
            pbe:LAPS_units="J/KG";

         //      negative buoyant energy         //

         float
            nbe(record,z,y,x);
            nbe:navigation_dim = "nav";
            nbe:record = "valtime, reftime";
            nbe:_FillValue = 1.e+37f;
            nbe:long_name="negative buoyant energy";
            nbe:units="joules/kilogram";
            nbe:valid_range= -20000.f, 20000.f;
            nbe:LAPS_var="NBE";
            nbe:lvl_coord="AGL";
            nbe:LAPS_units="J/KG";

        //      surface pressure        //

        float
            ps(record,z,y,x);
            ps:navigation_dim = "nav";
            ps:record = "valtime, reftime";
            ps:_FillValue = 1.e+37f;
            ps:long_name="surface pressure";
            ps:units="pascals";
            ps:valid_range= -20000.f, 20000.f;
            ps:LAPS_var="PS";
            ps:lvl_coord="AGL";
            ps:LAPS_units="PA";

        //      Cloud Ceiling           //

        float
            cce(record,z,y,x);
            cce:navigation_dim = "nav";
            cce:record = "valtime, reftime";
            cce:_FillValue = 1.e+37f;
            cce:long_name="cloud ceiling";
            cce:units="meters";
            cce:valid_range= -20000.f, 20000.f;
            cce:LAPS_var="CCE";
            cce:lvl_coord="AGL";
            cce:LAPS_units="M";

         //      visability              //

         float
            vis(record,z,y,x);
            vis:navigation_dim = "nav";
            vis:record = "valtime, reftime";
            vis:_FillValue = 1.e+37f;
            vis:long_name="visibility";
            vis:units="meters";
            vis:valid_range= -20000.f, 20000.f;
            vis:LAPS_var="VIS";
            vis:lvl_coord="AGL";
            vis:LAPS_units="M";

        //      LAPS cloud cover

        float
            lcv(record,z,y,x);
            lcv:navigation_dim = "nav";
            lcv:record = "valtime, reftime";
            lcv:_FillValue = 1.e+37f;
            lcv:long_name="LAPS cloud cover";
            lcv:units="none";
            lcv:valid_range= 0.f, 100.f;
            lcv:LAPS_var="LCV";
            lcv:lvl_coord="MSL";
            lcv:LAPS_units="UNDIM";

        //       Max echo tops

        float
            lmt(record,z,y,x);
            lmt:navigation_dim = "nav";
            lmt:record = "valtime, reftime";
            lmt:_FillValue = 1.e+37f;
            lmt:long_name="maximum radar echo tops";
            lmt:units="meters";
            lmt:valid_range= 0.f, 0.100f;
            lmt:LAPS_var="LMT";
            lmt:lvl_coord="MSL";
            lmt:LAPS_units="M";

        //      LAPS Fcst sfc precip type  //

        float
            spt(record,z,y,x);
            spt:navigation_dim = "nav";
            spt:record = "valtime, reftime";
            spt:_FillValue = 1.e+37f;
            spt:long_name="LAPS Fcst sfc precip type";
            spt:units="meters";
            spt:valid_range= 0.f, 0.100f;
            spt:LAPS_var="SPT";
            spt:lvl_coord="MSL";
            spt:LAPS_units="M";

        //      helicity

        float
            lhe(record,z,y,x);
            lhe:navigation_dim = "nav";
            lhe:record = "valtime, reftime";
            lhe:_FillValue = 1.e+37f;
            lhe:long_name="helicity";
            lhe:units="meters / second**2";
            lhe:valid_range= 0.f, 0.100f;
            lhe:LAPS_var="LHE";
            lhe:lvl_coord="MSL ";
            lhe:LAPS_units="M/S**2";

        //     lifted index            / 

        float
            li(record,z,y,x);
            li:navigation_dim = "nav";
            li:record = "valtime, reftime";
            li:_FillValue = 1.e+37f;
            li:long_name="lifted index";
            li:units="degrees Kelvin";
            li:valid_range= -20000.f, 20000.f;
            li:LAPS_var="LI";
            li:lvl_coord="AGL";
            li:LAPS_units="K";


         //      heat index                      //
         float
            hi(record,z,y,x);
            hi:navigation_dim = "nav";
            hi:record = "valtime, reftime";
            hi:_FillValue = 1.e+37f;
            hi:long_name="Heat index";
            hi:units="none";
            hi:valid_range= 0.f, 20.f;
            hi:LAPS_var="HI";
            hi:lvl_coord="none";
            hi:LAPS_units="none";

        //	LAPS variables
                	        
        long
            imax,
            jmax,
            kmax,
            kdim;

        char
            u_comment(record,z,namelen),
            v_comment(record,z,namelen),
            t_comment(record,z,namelen),
            p_comment(record,z,namelen),
            td_comment(record,z,namelen),
            rh_comment(record,z,namelen),
            lcb_comment(record,z,namelen),
            lct_comment(record,z,namelen),
            msl_comment(record,z,namelen),
            lil_comment(record,z,namelen),
            tpw_comment(record,z,namelen),
            r01_comment(record,z,namelen),
            rto_comment(record,z,namelen),
            s01_comment(record,z,namelen),
            sto_comment(record,z,namelen),
            th_comment(record,z,namelen),
            the_comment(record,z,namelen),
            pbe_comment(record,z,namelen),
            nbe_comment(record,z,namelen),
            ps_comment(record,z,namelen),
            cce_comment(record,z,namelen),
            vis_comment(record,z,namelen),
            lcv_comment(record,z,namelen),
            lmt_comment(record,z,namelen),
            spt_comment(record,z,namelen),
            lhe_comment(record,z,namelen),
            li_comment(record,z,namelen),
            hi_comment(record,z,namelen),
            asctime(record,namelen);

			
        //	inventory variables

        short
            u_fcinv(record, z);
            u_fcinv:_FillValue= 0s;
              	
        short
            v_fcinv(record, z);
            v_fcinv:_FillValue= 0s;
              	
        short
            p_fcinv(record, z);
            p_fcinv:_FillValue= 0s;
              	
        short
            t_fcinv(record, z);
            t_fcinv:_FillValue= 0s;
              	
        short
            td_fcinv(record, z);
            td_fcinv:_FillValue= 0s;
              	
        short
            rh_fcinv(record, z);
            rh_fcinv:_FillValue= 0s;

        short
            lcb_fcinv(record, z);
            lcb_fcinv:_FillValue= 0s;

        short
            lct_fcinv(record, z);
            lct_fcinv:_FillValue= 0s;

        short
            msl_fcinv(record, z);
            msl_fcinv:_FillValue= 0s;

        short
            lil_fcinv(record, z);
            lil_fcinv:_FillValue= 0s;

        short
            tpw_fcinv(record, z);
            tpw_fcinv:_FillValue= 0s;

        short
            r01_fcinv(record, z);
            r01_fcinv:_FillValue= 0s;

        short
            rto_fcinv(record, z);
            rto_fcinv:_FillValue= 0s;

        short
            s01_fcinv(record, z);
            s01_fcinv:_FillValue= 0s;

        short
            sto_fcinv(record, z);
            sto_fcinv:_FillValue= 0s;


        short
            th_fcinv(record, z);
            th_fcinv:_FillValue= 0s;

        short
            the_fcinv(record, z);
            the_fcinv:_FillValue= 0s;

        short
            pbe_fcinv(record, z);
            pbe_fcinv:_FillValue= 0s;

        short
            nbe_fcinv(record, z);
            nbe_fcinv:_FillValue= 0s;

        short
            ps_fcinv(record, z);
            ps_fcinv:_FillValue= 0s;

        short
            cce_fcinv(record, z);
            cce_fcinv:_FillValue= 0s;

        short
            vis_fcinv(record, z);
            vis_fcinv:_FillValue= 0s;

        short
            lcv_fcinv(record, z);
            lcv_fcinv:_FillValue= 0s;

        short
            lmt_fcinv(record, z);
            lmt_fcinv:_FillValue= 0s;

        short
            spt_fcinv(record, z);
            spt_fcinv:_FillValue= 0s;

        short
            lhe_fcinv(record, z);
            lhe_fcinv:_FillValue= 0s;

        short
            li_fcinv(record, z);
            li_fcinv:_FillValue= 0s;

        short
            hi_fcinv(record, z);
            hi_fcinv:_FillValue= 0s;


        //	list of grid levels

        float 
            level(z);
            level:long_name="level of data";
	    level:units = "hectopascals";
                    	
        //      validtime of the grid 

        double
            valtime(record);
            valtime:long_name = "valid time";
            valtime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      reference time of the process

        double
            reftime(record);
            reftime:long_name = "reference time";
            reftime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      nice name for originating center

        char
            origin_name(namelen);

        //      nice name for process

        char
            process_name(namelen);

        //      nice name for grid description instance
        char
            grid_name(namelen);

        //      basic assumption about earth shape
        char
            earth_shape(namelen);

        // navigation variables using 
        // WMO FM 92-VIII Ext.GRIB specification names
  
        char    grid_type(nav, namelen);
                grid_type:long_name = "GRIB-1 grid type";
  
        char    x_dim(nav, namelen);
                x_dim:long_name = "longitude dimension";
  
        char    y_dim(nav, namelen);
                y_dim:long_name = "latitude dimension";
  
        short   Nx(nav);
                Nx:long_name = "number of x points";
  
        short   Ny(nav);
                Ny:long_name =  "number of y points";
  
        float   La1(nav);
                La1:long_name = "first latitude";
                La1:units = "degrees_north";
  
        float   Lo1(nav);
                Lo1:long_name = "first longitude";
                Lo1:units = "degrees_east" ;
    
        float   LoV(nav);
                LoV:long_name = "orientation of grid" ;
                LoV:units = "degrees_east";
  
        float   Latin1(nav);
                Latin1:long_name = "orientation of grid" ;
                Latin1:units = "degrees_north";

        float   Latin2(nav);
                Latin2:long_name = "orientation of grid" ;
                Latin2:units = "degrees_north";

        float   Dx(nav);
                Dx:long_name = "x grid increment";
                Dx:units = "kilometers";
  
        float   Dy(nav);
                Dy:long_name = "y grid increment";
                Dy:units = "kilometers";
  
        // end of navigation variables

        :Conventions = "NUWG";
        :history = "created by LAPS Branch of FSL";
        :record = "valtime, reftime";
        :title = "RAMS rsf file - surface data";
        :version = 3;

    data:

        earth_shape     = "spherical radius";
        grid_name       = "RAMS rsf file - surface data";
        process_name    = "RAMS - Regional Atmospheric Modeling System";
        x_dim           = "x";
        y_dim           = "y";
}                       
