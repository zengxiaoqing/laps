netcdf lfr {

    dimensions:
        record = unlimited,
        z = 1,
	x = 249,
	y = 209,
        nav = 1,
        namelen = 132;
		
    variables:
        //	ventilation index

	float                                  
            vnt(record,z,y,x);
            vnt:navigation_dim = "nav";
            vnt:record = "valtime, reftime";
            vnt:_FillValue = 1.e+37f;
            vnt:long_name="ventilation index";
            vnt:units="meters**2 / second";
            vnt:valid_range= 0.f, 100000.f;
            vnt:LAPS_var="VNT";
            vnt:lvl_coord="NONE";
	    vnt:LAPS_units="M**2/S";
                	        
        //	boundary layer mean u component

	float                                  
            upb(record,z,y,x);
            upb:navigation_dim = "nav";
            upb:record = "valtime, reftime";
            upb:_FillValue = 1.e+37f;
            upb:long_name="boundary layer mean u component";
            upb:units="meters / second";
            upb:valid_range= -200.f, 200.f;
            upb:LAPS_var="UPB";
            upb:lvl_coord="NONE";
	    upb:LAPS_units="M/S";
                	        
        //	boundary layer mean v component

	float                                  
            vpb(record,z,y,x);
            vpb:navigation_dim = "nav";
            vpb:record = "valtime, reftime";
            vpb:_FillValue = 1.e+37f;
            vpb:long_name="boundary layer mean v component";
            vpb:units="meters / second";
            vpb:valid_range= -200.f, 200.f;
            vpb:LAPS_var="VPB";
            vpb:lvl_coord="NONE";
	    vpb:LAPS_units="M/S";
                	        
        //	mid-level haines index
        float 
            ham(record,z,y,x) ;
            ham:navigation_dim = "nav";
            ham:record = "valtime, reftime";
            ham:_FillValue = 1.e+37f;
            ham:long_name = "mid-level haines index" ;
            ham:units = "none" ;
            ham:valid_range = 0.f, 6.0f ;
            ham:LAPS_var = "HAM" ;
            ham:lvl_coord = "NONE" ;
            ham:LAPS_units = "NONE" ;
                	        
        //	high-level haines index
        float 
            hah(record,z,y,x) ;
            hah:navigation_dim = "nav";
            hah:record = "valtime, reftime";
            hah:_FillValue = 1.e+37f;
            hah:long_name = "high-level haines index" ;
            hah:units = "none" ;
            hah:valid_range = 0.f, 6.0f ;
            hah:LAPS_var = "HAH" ;
            hah:lvl_coord = "NONE" ;
            hah:LAPS_units = "NONE" ;

        //	Fosberg fire weather index
        float 
            fwi(record,z,y,x) ;
            fwi:navigation_dim = "nav";
            fwi:record = "valtime, reftime";
            fwi:_FillValue = 1.e+37f;
            fwi:long_name = "Fosberg Index" ;
            fwi:units = "none" ;
            fwi:valid_range = 0.f, 40.0f ;
            fwi:LAPS_var = "FWI" ;
            fwi:lvl_coord = "NONE" ;
            fwi:LAPS_units = "NONE" ;

        //	Critical fire weather index
        float 
            cwi(record,z,y,x) ;
            cwi:navigation_dim = "nav";
            cwi:record = "valtime, reftime";
            cwi:_FillValue = 1.e+37f;
            cwi:long_name = "critical fire weather index" ;
            cwi:units = "none" ;
            cwi:valid_range = 0.f, 1.0f ;
            cwi:LAPS_var = "CWI" ;
            cwi:lvl_coord = "NONE" ;
            cwi:LAPS_units = "NONE" ;

        //	LAPS variables

        long
            imax,
            jmax,
            kmax,
            kdim;

        char
            vnt_comment(record,z,namelen),
            upb_comment(record,z,namelen),
            vpb_comment(record,z,namelen),
            ham_comment(record,z,namelen),
            hah_comment(record,z,namelen),
            fwi_comment(record,z,namelen),
            cwi_comment(record,z,namelen),
            asctime(record,namelen);

			
        //	inventory variables

        short
            vnt_fcinv(record, z);
            vnt_fcinv:_FillValue= 0s;
              	
        short
            upb_fcinv(record, z);
            upb_fcinv:_FillValue= 0s;
              	
        short
            vpb_fcinv(record, z);
            vpb_fcinv:_FillValue= 0s;
              	
        short
            ham_fcinv(record, z);
            ham_fcinv:_FillValue= 0s;
              	
        short
            hah_fcinv(record, z);
            hah_fcinv:_FillValue= 0s;
              	
        short
            fwi_fcinv(record, z);
            fwi_fcinv:_FillValue= 0s;
              	
        short
            cwi_fcinv(record, z);
            cwi_fcinv:_FillValue= 0s;
              	
        //	list of grid levels

        float 
            level(z);
            level:long_name="level of data";
	    level:units = "none";
                    	
        //      validtime of the grid 

        double
            valtime(record);
            valtime:long_name = "valid time";
            valtime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      reference time of the process

        double
            reftime(record);
            reftime:long_name = "reference time";
            reftime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      nice name for originating center

        char
            origin_name(namelen);

        //      nice name for process

        char
            process_name(namelen);

        //      nice name for grid description instance
        char
            grid_name(namelen);

        //      basic assumption about earth shape
        char
            earth_shape(namelen);

        // navigation variables using 
        // WMO FM 92-VIII Ext.GRIB specification names
  
        char    grid_type(nav, namelen);
                grid_type:long_name = "GRIB-1 grid type";
  
        char    x_dim(nav, namelen);
                x_dim:long_name = "longitude dimension";
  
        char    y_dim(nav, namelen);
                y_dim:long_name = "latitude dimension";
  
        short   Nx(nav);
                Nx:long_name = "number of x points";
  
        short   Ny(nav);
                Ny:long_name =  "number of y points";
  
        float   La1(nav);
                La1:long_name = "first latitude";
                La1:units = "degrees_north";
  
        float   Lo1(nav);
                Lo1:long_name = "first longitude";
                Lo1:units = "degrees_east" ;
    
        float   LoV(nav);
                LoV:long_name = "orientation of grid" ;
                LoV:units = "degrees_east";
  
        float   Latin1(nav);
                Latin1:long_name = "orientation of grid" ;
                Latin1:units = "degrees_north";

        float   Latin2(nav);
                Latin2:long_name = "orientation of grid" ;
                Latin2:units = "degrees_north";

        float   Dx(nav);
                Dx:long_name = "x grid increment";
                Dx:units = "meters";
  
        float   Dy(nav);
                Dy:long_name = "y grid increment";
                Dy:units = "meters";
  
        // end of navigation variables

        :Conventions = "NUWG";
        :history = "created by LAPS Branch of FSL";
        :record = "valtime, reftime";
        :title = "LAPS lfr file - fire weather";
        :version = 3;

    data:

        earth_shape     = "spherical radius";
        grid_name       = "LAPS lfr file - fire weather";
        process_name    = "LAPS - Local Analysis and Prediction System";
        x_dim           = "x";
        y_dim           = "y";
}                       
